module CHIP(    
	// Input signals
    clk,
    rst_n,
	in_valid,
    in_valid_num,
    col,
    row,
    in_num,
	
    // Output signals
	out_valid,
    out
);

// ===============================================================
// Input & Output Declaration
// ===============================================================
input           clk, rst_n, in_valid,in_valid_num;
input   [3:0]   col,row;
input   [2:0]   in_num;

output          out_valid;
output  [3:0]   out;

wire		    C_clk;
wire			C_rst_n;
wire			C_in_valid;
wire			C_in_valid_num;
wire	[3:0]	C_col;
wire	[3:0]	C_row;
wire	[2:0]	C_in_num;

wire			C_out_valid;
wire	[3:0]	C_out;


wire	        BUF_clk;
CLKBUFX20 buf0(.A(C_clk),.Y(BUF_clk));


QUEEN u_QUEEN(
    .clk(BUF_clk),
    .rst_n(C_rst_n),
    .in_valid(C_in_valid),
    .in_valid_num(C_in_valid_num),
    .col(C_col),
    .row(C_row),
    .in_num(C_in_num),

    .out_valid(C_out_valid),
    .out(C_out)
);

//////////////
P8C I_CLK      ( .Y(C_clk),        .P(clk),        .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b0), .CSEN(1'b1) );
P8C I_RESET    ( .Y(C_rst_n),      .P(rst_n),      .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_IN_VALID    ( .Y(C_in_valid),   .P(in_valid),   .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_IN_VALID_NUM    ( .Y(C_in_valid_num),   .P(in_valid_num),   .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_COL_0     ( .Y(C_col[0]), .P(col[0]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_COL_1     ( .Y(C_col[1]), .P(col[1]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_COL_2     ( .Y(C_col[2]), .P(col[2]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_COL_3     ( .Y(C_col[3]), .P(col[3]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_ROW_0     ( .Y(C_row[0]), .P(row[0]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_ROW_1     ( .Y(C_row[1]), .P(row[1]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_ROW_2     ( .Y(C_row[2]), .P(row[2]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_ROW_3     ( .Y(C_row[3]), .P(row[3]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_IN_NUM_0     ( .Y(C_in_num[0]), .P(in_num[0]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_IN_NUM_1     ( .Y(C_in_num[1]), .P(in_num[1]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_IN_NUM_2     ( .Y(C_in_num[2]), .P(in_num[2]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );

P8C O_OUT_VALID    ( .A(C_out_valid), 	.P(out_valid), 	 .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0));
P8C O_OUT_0     ( .A(C_out[0]),   	.P(out[0]), 	.ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0));
P8C O_OUT_1     ( .A(C_out[1]),   	.P(out[1]), 	.ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0));
P8C O_OUT_2     ( .A(C_out[2]),   	.P(out[2]), 	.ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0));
P8C O_OUT_3     ( .A(C_out[3]),   	.P(out[3]), 	.ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0));



//I/O power 3.3V pads x8 (DVDD + DGND)
PVDDR VDDP0 ();
PVSSR GNDP0 ();
PVDDR VDDP1 ();
PVSSR GNDP1 ();
PVDDR VDDP2 ();
PVSSR GNDP2 ();
PVDDR VDDP3 ();
PVSSR GNDP3 ();
PVDDR VDDP4 ();
PVSSR GNDP4 ();
PVDDR VDDP5 ();
PVSSR GNDP5 ();
PVDDR VDDP6 ();
PVSSR GNDP6 ();
PVDDR VDDP7 ();
PVSSR GNDP7 ();

//Core poweri 1.8V pads x8 (VDD + GND)
PVDDC VDDC0 ();
PVSSC GNDC0 ();
PVDDC VDDC1 ();
PVSSC GNDC1 ();
PVDDC VDDC2 ();
PVSSC GNDC2 ();
PVDDC VDDC3 ();
PVSSC GNDC3 ();
PVDDC VDDC4 ();
PVSSC GNDC4 ();
PVDDC VDDC5 ();
PVSSC GNDC5 ();
PVDDC VDDC6 ();
PVSSC GNDC6 ();
PVDDC VDDC7 ();
PVSSC GNDC7 ();


endmodule/////////////////////////////////////////////////////////////
// Created by: Synopsys DC Ultra(TM) in wire load mode
// Version   : T-2022.03
// Date      : Thu May  4 22:05:21 2023
/////////////////////////////////////////////////////////////


module QUEEN ( clk, rst_n, in_valid, col, row, in_valid_num, in_num, out_valid, 
        out, Port10 );
  input [3:0] col;
  input [3:0] row;
  input [2:0] in_num;
  output [3:0] out;
  input clk, rst_n, in_valid, in_valid_num, Port10;
  output out_valid;
  wire   N4586, N6082, N6083, N6084, N6085, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
         n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
         n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
         n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
         n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
         n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
         n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
         n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
         n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
         n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
         n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
         n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
         n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
         n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
         n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
         n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
         n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
         n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
         n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
         n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
         n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
         n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
         n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
         n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
         n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
         n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
         n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
         n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086;
  wire   [2:0] current_state;
  wire   [3:0] count_receive;
  wire   [3:1] count;
  wire   [3:0] count_out;
  wire   [2:0] x;
  wire   [11:0] array_in;
  wire   [47:0] row_store;
  wire   [11:0] x_array;
  wire   [11:0] y_array;
  wire   [22:0] sub_array;
  wire   [22:0] add_array;
  wire   [143:0] array_look_back;

  DFFRHQXL count_out_reg_1_ ( .D(N6083), .CK(clk), .RN(rst_n), .Q(count_out[1]) );
  DFFRHQXL count_out_reg_2_ ( .D(N6084), .CK(clk), .RN(rst_n), .Q(count_out[2]) );
  DFFRHQXL current_state_reg_2_ ( .D(n1683), .CK(clk), .RN(rst_n), .Q(
        current_state[2]) );
  DFFRHQXL count_receive_reg_0_ ( .D(n1679), .CK(clk), .RN(rst_n), .Q(
        count_receive[0]) );
  DFFRHQXL count_receive_reg_1_ ( .D(n1678), .CK(clk), .RN(rst_n), .Q(
        count_receive[1]) );
  DFFRHQXL count_receive_reg_2_ ( .D(n1677), .CK(clk), .RN(rst_n), .Q(
        count_receive[2]) );
  DFFRHQXL count_receive_reg_3_ ( .D(n1676), .CK(clk), .RN(rst_n), .Q(
        count_receive[3]) );
  DFFRHQXL array_in_reg_0_ ( .D(n1675), .CK(clk), .RN(rst_n), .Q(array_in[0])
         );
  DFFRHQXL array_in_reg_2_ ( .D(n1673), .CK(clk), .RN(rst_n), .Q(array_in[2])
         );
  DFFRHQXL array_in_reg_3_ ( .D(n1672), .CK(clk), .RN(rst_n), .Q(array_in[3])
         );
  DFFRHQXL array_in_reg_4_ ( .D(n1671), .CK(clk), .RN(rst_n), .Q(array_in[4])
         );
  DFFRHQXL array_in_reg_5_ ( .D(n1670), .CK(clk), .RN(rst_n), .Q(array_in[5])
         );
  DFFRHQXL array_in_reg_6_ ( .D(n1669), .CK(clk), .RN(rst_n), .Q(array_in[6])
         );
  DFFRHQXL array_in_reg_7_ ( .D(n1668), .CK(clk), .RN(rst_n), .Q(array_in[7])
         );
  DFFRHQXL array_in_reg_8_ ( .D(n1667), .CK(clk), .RN(rst_n), .Q(array_in[8])
         );
  DFFRHQXL array_in_reg_9_ ( .D(n1666), .CK(clk), .RN(rst_n), .Q(array_in[9])
         );
  DFFRHQXL array_in_reg_10_ ( .D(n1665), .CK(clk), .RN(rst_n), .Q(array_in[10]) );
  DFFRHQXL array_in_reg_11_ ( .D(n1664), .CK(clk), .RN(rst_n), .Q(array_in[11]) );
  DFFRHQXL array_in_reg_1_ ( .D(n1674), .CK(clk), .RN(rst_n), .Q(array_in[1])
         );
  DFFRHQXL y_array_reg_4_ ( .D(n1400), .CK(clk), .RN(rst_n), .Q(y_array[4]) );
  DFFRHQX4 x_reg_0_ ( .D(n1613), .CK(clk), .RN(rst_n), .Q(x[0]) );
  DFFRHQX4 x_reg_1_ ( .D(n1614), .CK(clk), .RN(rst_n), .Q(x[1]) );
  DFFRHQXL current_state_reg_1_ ( .D(n1684), .CK(clk), .RN(rst_n), .Q(
        current_state[1]) );
  DFFRHQXL current_state_reg_0_ ( .D(n1685), .CK(clk), .RN(rst_n), .Q(
        current_state[0]) );
  DFFRHQXL row_store_reg_10__1_ ( .D(n1620), .CK(clk), .RN(rst_n), .Q(
        row_store[41]) );
  DFFRHQXL row_store_reg_8__1_ ( .D(n1628), .CK(clk), .RN(rst_n), .Q(
        row_store[33]) );
  DFFRHQXL row_store_reg_7__1_ ( .D(n1632), .CK(clk), .RN(rst_n), .Q(
        row_store[29]) );
  DFFRHQXL row_store_reg_5__1_ ( .D(n1640), .CK(clk), .RN(rst_n), .Q(
        row_store[21]) );
  DFFRHQXL row_store_reg_4__1_ ( .D(n1644), .CK(clk), .RN(rst_n), .Q(
        row_store[17]) );
  DFFRHQXL row_store_reg_6__1_ ( .D(n1636), .CK(clk), .RN(rst_n), .Q(
        row_store[25]) );
  DFFRHQXL row_store_reg_2__1_ ( .D(n1652), .CK(clk), .RN(rst_n), .Q(
        row_store[9]) );
  DFFRHQXL row_store_reg_11__1_ ( .D(n1616), .CK(clk), .RN(rst_n), .Q(
        row_store[45]) );
  DFFRHQXL row_store_reg_9__1_ ( .D(n1624), .CK(clk), .RN(rst_n), .Q(
        row_store[37]) );
  DFFRHQXL row_store_reg_3__1_ ( .D(n1648), .CK(clk), .RN(rst_n), .Q(
        row_store[13]) );
  DFFRHQXL row_store_reg_1__1_ ( .D(n1656), .CK(clk), .RN(rst_n), .Q(
        row_store[5]) );
  DFFRHQXL row_store_reg_1__3_ ( .D(n1658), .CK(clk), .RN(rst_n), .Q(
        row_store[7]) );
  DFFRHQXL row_store_reg_2__3_ ( .D(n1654), .CK(clk), .RN(rst_n), .Q(
        row_store[11]) );
  DFFRHQXL row_store_reg_3__3_ ( .D(n1650), .CK(clk), .RN(rst_n), .Q(
        row_store[15]) );
  DFFRHQXL row_store_reg_4__3_ ( .D(n1646), .CK(clk), .RN(rst_n), .Q(
        row_store[19]) );
  DFFRHQXL row_store_reg_5__3_ ( .D(n1642), .CK(clk), .RN(rst_n), .Q(
        row_store[23]) );
  DFFRHQXL row_store_reg_6__3_ ( .D(n1638), .CK(clk), .RN(rst_n), .Q(
        row_store[27]) );
  DFFRHQXL row_store_reg_7__3_ ( .D(n1634), .CK(clk), .RN(rst_n), .Q(
        row_store[31]) );
  DFFRHQXL row_store_reg_8__3_ ( .D(n1630), .CK(clk), .RN(rst_n), .Q(
        row_store[35]) );
  DFFRHQXL row_store_reg_9__3_ ( .D(n1626), .CK(clk), .RN(rst_n), .Q(
        row_store[39]) );
  DFFRHQXL row_store_reg_10__3_ ( .D(n1622), .CK(clk), .RN(rst_n), .Q(
        row_store[43]) );
  DFFRHQXL row_store_reg_11__3_ ( .D(n1618), .CK(clk), .RN(rst_n), .Q(
        row_store[47]) );
  DFFRHQXL row_store_reg_1__0_ ( .D(n1659), .CK(clk), .RN(rst_n), .Q(
        row_store[4]) );
  DFFRHQXL row_store_reg_2__0_ ( .D(n1655), .CK(clk), .RN(rst_n), .Q(
        row_store[8]) );
  DFFRHQXL row_store_reg_3__0_ ( .D(n1651), .CK(clk), .RN(rst_n), .Q(
        row_store[12]) );
  DFFRHQXL row_store_reg_4__0_ ( .D(n1647), .CK(clk), .RN(rst_n), .Q(
        row_store[16]) );
  DFFRHQXL row_store_reg_5__0_ ( .D(n1643), .CK(clk), .RN(rst_n), .Q(
        row_store[20]) );
  DFFRHQXL row_store_reg_6__0_ ( .D(n1639), .CK(clk), .RN(rst_n), .Q(
        row_store[24]) );
  DFFRHQXL row_store_reg_7__0_ ( .D(n1635), .CK(clk), .RN(rst_n), .Q(
        row_store[28]) );
  DFFRHQXL row_store_reg_8__0_ ( .D(n1631), .CK(clk), .RN(rst_n), .Q(
        row_store[32]) );
  DFFRHQXL row_store_reg_9__0_ ( .D(n1627), .CK(clk), .RN(rst_n), .Q(
        row_store[36]) );
  DFFRHQXL row_store_reg_10__0_ ( .D(n1623), .CK(clk), .RN(rst_n), .Q(
        row_store[40]) );
  DFFRHQXL row_store_reg_11__0_ ( .D(n1619), .CK(clk), .RN(rst_n), .Q(
        row_store[44]) );
  DFFRHQXL row_store_reg_1__2_ ( .D(n1657), .CK(clk), .RN(rst_n), .Q(
        row_store[6]) );
  DFFRHQXL row_store_reg_2__2_ ( .D(n1653), .CK(clk), .RN(rst_n), .Q(
        row_store[10]) );
  DFFRHQXL row_store_reg_3__2_ ( .D(n1649), .CK(clk), .RN(rst_n), .Q(
        row_store[14]) );
  DFFRHQXL row_store_reg_4__2_ ( .D(n1645), .CK(clk), .RN(rst_n), .Q(
        row_store[18]) );
  DFFRHQXL row_store_reg_5__2_ ( .D(n1641), .CK(clk), .RN(rst_n), .Q(
        row_store[22]) );
  DFFRHQXL row_store_reg_6__2_ ( .D(n1637), .CK(clk), .RN(rst_n), .Q(
        row_store[26]) );
  DFFRHQXL row_store_reg_7__2_ ( .D(n1633), .CK(clk), .RN(rst_n), .Q(
        row_store[30]) );
  DFFRHQXL row_store_reg_8__2_ ( .D(n1629), .CK(clk), .RN(rst_n), .Q(
        row_store[34]) );
  DFFRHQXL row_store_reg_9__2_ ( .D(n1625), .CK(clk), .RN(rst_n), .Q(
        row_store[38]) );
  DFFRHQXL row_store_reg_10__2_ ( .D(n1621), .CK(clk), .RN(rst_n), .Q(
        row_store[42]) );
  DFFRHQXL row_store_reg_11__2_ ( .D(n1617), .CK(clk), .RN(rst_n), .Q(
        row_store[46]) );
  DFFRHQXL x_array_reg_11_ ( .D(n1612), .CK(clk), .RN(rst_n), .Q(x_array[11])
         );
  DFFRHQXL x_array_reg_10_ ( .D(n1611), .CK(clk), .RN(rst_n), .Q(x_array[10])
         );
  DFFRHQXL x_array_reg_9_ ( .D(n1610), .CK(clk), .RN(rst_n), .Q(x_array[9]) );
  DFFRHQXL x_array_reg_8_ ( .D(n1609), .CK(clk), .RN(rst_n), .Q(x_array[8]) );
  DFFRHQXL x_array_reg_7_ ( .D(n1608), .CK(clk), .RN(rst_n), .Q(x_array[7]) );
  DFFRHQXL x_array_reg_6_ ( .D(n1607), .CK(clk), .RN(rst_n), .Q(x_array[6]) );
  DFFRHQXL x_array_reg_5_ ( .D(n1606), .CK(clk), .RN(rst_n), .Q(x_array[5]) );
  DFFRHQXL x_array_reg_4_ ( .D(n1605), .CK(clk), .RN(rst_n), .Q(x_array[4]) );
  DFFRHQXL x_array_reg_3_ ( .D(n1604), .CK(clk), .RN(rst_n), .Q(x_array[3]) );
  DFFRHQXL x_array_reg_2_ ( .D(n1603), .CK(clk), .RN(rst_n), .Q(x_array[2]) );
  DFFRHQXL x_array_reg_1_ ( .D(n1602), .CK(clk), .RN(rst_n), .Q(x_array[1]) );
  DFFRHQXL x_array_reg_0_ ( .D(n1601), .CK(clk), .RN(rst_n), .Q(x_array[0]) );
  DFFRHQXL sub_array_reg_11_ ( .D(n1453), .CK(clk), .RN(rst_n), .Q(
        sub_array[11]) );
  DFFRHQXL sub_array_reg_12_ ( .D(n1452), .CK(clk), .RN(rst_n), .Q(
        sub_array[12]) );
  DFFRHQXL sub_array_reg_13_ ( .D(n1451), .CK(clk), .RN(rst_n), .Q(
        sub_array[13]) );
  DFFRHQXL sub_array_reg_14_ ( .D(n1450), .CK(clk), .RN(rst_n), .Q(
        sub_array[14]) );
  DFFRHQXL sub_array_reg_15_ ( .D(n1449), .CK(clk), .RN(rst_n), .Q(
        sub_array[15]) );
  DFFRHQXL sub_array_reg_16_ ( .D(n1448), .CK(clk), .RN(rst_n), .Q(
        sub_array[16]) );
  DFFRHQXL sub_array_reg_17_ ( .D(n1447), .CK(clk), .RN(rst_n), .Q(
        sub_array[17]) );
  DFFRHQXL sub_array_reg_18_ ( .D(n1446), .CK(clk), .RN(rst_n), .Q(
        sub_array[18]) );
  DFFRHQXL sub_array_reg_19_ ( .D(n1445), .CK(clk), .RN(rst_n), .Q(
        sub_array[19]) );
  DFFRHQXL sub_array_reg_20_ ( .D(n1444), .CK(clk), .RN(rst_n), .Q(
        sub_array[20]) );
  DFFRHQXL sub_array_reg_21_ ( .D(n1443), .CK(clk), .RN(rst_n), .Q(
        sub_array[21]) );
  DFFRHQXL sub_array_reg_22_ ( .D(n1442), .CK(clk), .RN(rst_n), .Q(
        sub_array[22]) );
  DFFRHQXL sub_array_reg_3_ ( .D(n1441), .CK(clk), .RN(rst_n), .Q(sub_array[3]) );
  DFFRHQXL sub_array_reg_4_ ( .D(n1440), .CK(clk), .RN(rst_n), .Q(sub_array[4]) );
  DFFRHQXL sub_array_reg_5_ ( .D(n1439), .CK(clk), .RN(rst_n), .Q(sub_array[5]) );
  DFFRHQXL sub_array_reg_6_ ( .D(n1438), .CK(clk), .RN(rst_n), .Q(sub_array[6]) );
  DFFRHQXL sub_array_reg_7_ ( .D(n1437), .CK(clk), .RN(rst_n), .Q(sub_array[7]) );
  DFFRHQXL sub_array_reg_1_ ( .D(n1436), .CK(clk), .RN(rst_n), .Q(sub_array[1]) );
  DFFRHQXL sub_array_reg_9_ ( .D(n1435), .CK(clk), .RN(rst_n), .Q(sub_array[9]) );
  DFFRHQXL sub_array_reg_0_ ( .D(n1434), .CK(clk), .RN(rst_n), .Q(sub_array[0]) );
  DFFRHQXL sub_array_reg_2_ ( .D(n1433), .CK(clk), .RN(rst_n), .Q(sub_array[2]) );
  DFFRHQXL sub_array_reg_8_ ( .D(n1432), .CK(clk), .RN(rst_n), .Q(sub_array[8]) );
  DFFRHQXL sub_array_reg_10_ ( .D(n1431), .CK(clk), .RN(rst_n), .Q(
        sub_array[10]) );
  DFFRHQXL add_array_reg_0_ ( .D(n1430), .CK(clk), .RN(rst_n), .Q(add_array[0]) );
  DFFRHQXL add_array_reg_2_ ( .D(n1429), .CK(clk), .RN(rst_n), .Q(add_array[2]) );
  DFFRHQXL add_array_reg_4_ ( .D(n1428), .CK(clk), .RN(rst_n), .Q(add_array[4]) );
  DFFRHQXL add_array_reg_6_ ( .D(n1427), .CK(clk), .RN(rst_n), .Q(add_array[6]) );
  DFFRHQXL add_array_reg_8_ ( .D(n1426), .CK(clk), .RN(rst_n), .Q(add_array[8]) );
  DFFRHQXL add_array_reg_10_ ( .D(n1425), .CK(clk), .RN(rst_n), .Q(
        add_array[10]) );
  DFFRHQXL add_array_reg_12_ ( .D(n1424), .CK(clk), .RN(rst_n), .Q(
        add_array[12]) );
  DFFRHQXL add_array_reg_14_ ( .D(n1423), .CK(clk), .RN(rst_n), .Q(
        add_array[14]) );
  DFFRHQXL add_array_reg_1_ ( .D(n1422), .CK(clk), .RN(rst_n), .Q(add_array[1]) );
  DFFRHQXL add_array_reg_3_ ( .D(n1421), .CK(clk), .RN(rst_n), .Q(add_array[3]) );
  DFFRHQXL add_array_reg_5_ ( .D(n1420), .CK(clk), .RN(rst_n), .Q(add_array[5]) );
  DFFRHQXL add_array_reg_7_ ( .D(n1419), .CK(clk), .RN(rst_n), .Q(add_array[7]) );
  DFFRHQXL add_array_reg_9_ ( .D(n1418), .CK(clk), .RN(rst_n), .Q(add_array[9]) );
  DFFRHQXL add_array_reg_11_ ( .D(n1417), .CK(clk), .RN(rst_n), .Q(
        add_array[11]) );
  DFFRHQXL add_array_reg_13_ ( .D(n1416), .CK(clk), .RN(rst_n), .Q(
        add_array[13]) );
  DFFRHQXL add_array_reg_15_ ( .D(n1415), .CK(clk), .RN(rst_n), .Q(
        add_array[15]) );
  DFFRHQXL add_array_reg_17_ ( .D(n1414), .CK(clk), .RN(rst_n), .Q(
        add_array[17]) );
  DFFRHQXL add_array_reg_19_ ( .D(n1413), .CK(clk), .RN(rst_n), .Q(
        add_array[19]) );
  DFFRHQXL add_array_reg_21_ ( .D(n1412), .CK(clk), .RN(rst_n), .Q(
        add_array[21]) );
  DFFRHQXL add_array_reg_16_ ( .D(n1411), .CK(clk), .RN(rst_n), .Q(
        add_array[16]) );
  DFFRHQXL add_array_reg_18_ ( .D(n1410), .CK(clk), .RN(rst_n), .Q(
        add_array[18]) );
  DFFRHQXL add_array_reg_20_ ( .D(n1409), .CK(clk), .RN(rst_n), .Q(
        add_array[20]) );
  DFFRHQXL add_array_reg_22_ ( .D(n1408), .CK(clk), .RN(rst_n), .Q(
        add_array[22]) );
  DFFRHQXL y_array_reg_5_ ( .D(n1401), .CK(clk), .RN(rst_n), .Q(y_array[5]) );
  DFFRHQXL array_look_back_reg_0__4_ ( .D(n1469), .CK(clk), .RN(rst_n), .Q(
        array_look_back[4]) );
  DFFRHQXL array_look_back_reg_1__4_ ( .D(n1468), .CK(clk), .RN(rst_n), .Q(
        array_look_back[16]) );
  DFFRHQXL array_look_back_reg_2__4_ ( .D(n1467), .CK(clk), .RN(rst_n), .Q(
        array_look_back[28]) );
  DFFRHQXL array_look_back_reg_3__4_ ( .D(n1466), .CK(clk), .RN(rst_n), .Q(
        array_look_back[40]) );
  DFFRHQXL array_look_back_reg_4__4_ ( .D(n1465), .CK(clk), .RN(rst_n), .Q(
        array_look_back[52]) );
  DFFRHQXL array_look_back_reg_5__4_ ( .D(n1464), .CK(clk), .RN(rst_n), .Q(
        array_look_back[64]) );
  DFFRHQXL array_look_back_reg_6__4_ ( .D(n1463), .CK(clk), .RN(rst_n), .Q(
        array_look_back[76]) );
  DFFRHQXL array_look_back_reg_7__4_ ( .D(n1462), .CK(clk), .RN(rst_n), .Q(
        array_look_back[88]) );
  DFFRHQXL array_look_back_reg_8__4_ ( .D(n1461), .CK(clk), .RN(rst_n), .Q(
        array_look_back[100]) );
  DFFRHQXL array_look_back_reg_9__4_ ( .D(n1460), .CK(clk), .RN(rst_n), .Q(
        array_look_back[112]) );
  DFFRHQXL array_look_back_reg_10__4_ ( .D(n1459), .CK(clk), .RN(rst_n), .Q(
        array_look_back[124]) );
  DFFRHQXL array_look_back_reg_11__4_ ( .D(n1458), .CK(clk), .RN(rst_n), .Q(
        array_look_back[136]) );
  DFFRHQXL y_array_reg_0_ ( .D(n1404), .CK(clk), .RN(rst_n), .Q(y_array[0]) );
  DFFRHQXL array_look_back_reg_0__7_ ( .D(n1505), .CK(clk), .RN(rst_n), .Q(
        array_look_back[7]) );
  DFFRHQXL array_look_back_reg_1__7_ ( .D(n1504), .CK(clk), .RN(rst_n), .Q(
        array_look_back[19]) );
  DFFRHQXL array_look_back_reg_2__7_ ( .D(n1503), .CK(clk), .RN(rst_n), .Q(
        array_look_back[31]) );
  DFFRHQXL array_look_back_reg_3__7_ ( .D(n1502), .CK(clk), .RN(rst_n), .Q(
        array_look_back[43]) );
  DFFRHQXL array_look_back_reg_4__7_ ( .D(n1501), .CK(clk), .RN(rst_n), .Q(
        array_look_back[55]) );
  DFFRHQXL array_look_back_reg_5__7_ ( .D(n1500), .CK(clk), .RN(rst_n), .Q(
        array_look_back[67]) );
  DFFRHQXL array_look_back_reg_6__7_ ( .D(n1499), .CK(clk), .RN(rst_n), .Q(
        array_look_back[79]) );
  DFFRHQXL array_look_back_reg_7__7_ ( .D(n1498), .CK(clk), .RN(rst_n), .Q(
        array_look_back[91]) );
  DFFRHQXL array_look_back_reg_8__7_ ( .D(n1497), .CK(clk), .RN(rst_n), .Q(
        array_look_back[103]) );
  DFFRHQXL array_look_back_reg_9__7_ ( .D(n1496), .CK(clk), .RN(rst_n), .Q(
        array_look_back[115]) );
  DFFRHQXL array_look_back_reg_10__7_ ( .D(n1495), .CK(clk), .RN(rst_n), .Q(
        array_look_back[127]) );
  DFFRHQXL array_look_back_reg_11__7_ ( .D(n1494), .CK(clk), .RN(rst_n), .Q(
        array_look_back[139]) );
  DFFRHQXL y_array_reg_7_ ( .D(n1403), .CK(clk), .RN(rst_n), .Q(y_array[7]) );
  DFFRHQXL array_look_back_reg_0__9_ ( .D(n1599), .CK(clk), .RN(rst_n), .Q(
        array_look_back[9]) );
  DFFRHQXL array_look_back_reg_1__9_ ( .D(n1595), .CK(clk), .RN(rst_n), .Q(
        array_look_back[21]) );
  DFFRHQXL array_look_back_reg_2__9_ ( .D(n1591), .CK(clk), .RN(rst_n), .Q(
        array_look_back[33]) );
  DFFRHQXL array_look_back_reg_3__9_ ( .D(n1587), .CK(clk), .RN(rst_n), .Q(
        array_look_back[45]) );
  DFFRHQXL array_look_back_reg_4__9_ ( .D(n1583), .CK(clk), .RN(rst_n), .Q(
        array_look_back[57]) );
  DFFRHQXL array_look_back_reg_5__9_ ( .D(n1579), .CK(clk), .RN(rst_n), .Q(
        array_look_back[69]) );
  DFFRHQXL array_look_back_reg_6__9_ ( .D(n1575), .CK(clk), .RN(rst_n), .Q(
        array_look_back[81]) );
  DFFRHQXL array_look_back_reg_7__9_ ( .D(n1571), .CK(clk), .RN(rst_n), .Q(
        array_look_back[93]) );
  DFFRHQXL array_look_back_reg_8__9_ ( .D(n1567), .CK(clk), .RN(rst_n), .Q(
        array_look_back[105]) );
  DFFRHQXL array_look_back_reg_9__9_ ( .D(n1563), .CK(clk), .RN(rst_n), .Q(
        array_look_back[117]) );
  DFFRHQXL array_look_back_reg_10__9_ ( .D(n1559), .CK(clk), .RN(rst_n), .Q(
        array_look_back[129]) );
  DFFRHQXL array_look_back_reg_11__9_ ( .D(n1555), .CK(clk), .RN(rst_n), .Q(
        array_look_back[141]) );
  DFFRHQXL array_look_back_reg_0__8_ ( .D(n1600), .CK(clk), .RN(rst_n), .Q(
        array_look_back[8]) );
  DFFRHQXL array_look_back_reg_1__8_ ( .D(n1596), .CK(clk), .RN(rst_n), .Q(
        array_look_back[20]) );
  DFFRHQXL array_look_back_reg_2__8_ ( .D(n1592), .CK(clk), .RN(rst_n), .Q(
        array_look_back[32]) );
  DFFRHQXL array_look_back_reg_3__8_ ( .D(n1588), .CK(clk), .RN(rst_n), .Q(
        array_look_back[44]) );
  DFFRHQXL array_look_back_reg_4__8_ ( .D(n1584), .CK(clk), .RN(rst_n), .Q(
        array_look_back[56]) );
  DFFRHQXL array_look_back_reg_5__8_ ( .D(n1580), .CK(clk), .RN(rst_n), .Q(
        array_look_back[68]) );
  DFFRHQXL array_look_back_reg_6__8_ ( .D(n1576), .CK(clk), .RN(rst_n), .Q(
        array_look_back[80]) );
  DFFRHQXL array_look_back_reg_7__8_ ( .D(n1572), .CK(clk), .RN(rst_n), .Q(
        array_look_back[92]) );
  DFFRHQXL array_look_back_reg_8__8_ ( .D(n1568), .CK(clk), .RN(rst_n), .Q(
        array_look_back[104]) );
  DFFRHQXL array_look_back_reg_9__8_ ( .D(n1564), .CK(clk), .RN(rst_n), .Q(
        array_look_back[116]) );
  DFFRHQXL array_look_back_reg_10__8_ ( .D(n1560), .CK(clk), .RN(rst_n), .Q(
        array_look_back[128]) );
  DFFRHQXL array_look_back_reg_11__8_ ( .D(n1556), .CK(clk), .RN(rst_n), .Q(
        array_look_back[140]) );
  DFFRHQXL array_look_back_reg_0__10_ ( .D(n1598), .CK(clk), .RN(rst_n), .Q(
        array_look_back[10]) );
  DFFRHQXL array_look_back_reg_1__10_ ( .D(n1594), .CK(clk), .RN(rst_n), .Q(
        array_look_back[22]) );
  DFFRHQXL array_look_back_reg_2__10_ ( .D(n1590), .CK(clk), .RN(rst_n), .Q(
        array_look_back[34]) );
  DFFRHQXL array_look_back_reg_3__10_ ( .D(n1586), .CK(clk), .RN(rst_n), .Q(
        array_look_back[46]) );
  DFFRHQXL array_look_back_reg_4__10_ ( .D(n1582), .CK(clk), .RN(rst_n), .Q(
        array_look_back[58]) );
  DFFRHQXL array_look_back_reg_5__10_ ( .D(n1578), .CK(clk), .RN(rst_n), .Q(
        array_look_back[70]) );
  DFFRHQXL array_look_back_reg_6__10_ ( .D(n1574), .CK(clk), .RN(rst_n), .Q(
        array_look_back[82]) );
  DFFRHQXL array_look_back_reg_7__10_ ( .D(n1570), .CK(clk), .RN(rst_n), .Q(
        array_look_back[94]) );
  DFFRHQXL array_look_back_reg_8__10_ ( .D(n1566), .CK(clk), .RN(rst_n), .Q(
        array_look_back[106]) );
  DFFRHQXL array_look_back_reg_9__10_ ( .D(n1562), .CK(clk), .RN(rst_n), .Q(
        array_look_back[118]) );
  DFFRHQXL array_look_back_reg_10__10_ ( .D(n1558), .CK(clk), .RN(rst_n), .Q(
        array_look_back[130]) );
  DFFRHQXL array_look_back_reg_11__10_ ( .D(n1554), .CK(clk), .RN(rst_n), .Q(
        array_look_back[142]) );
  DFFRHQXL array_look_back_reg_0__2_ ( .D(n1541), .CK(clk), .RN(rst_n), .Q(
        array_look_back[2]) );
  DFFRHQXL array_look_back_reg_1__2_ ( .D(n1540), .CK(clk), .RN(rst_n), .Q(
        array_look_back[14]) );
  DFFRHQXL array_look_back_reg_2__2_ ( .D(n1539), .CK(clk), .RN(rst_n), .Q(
        array_look_back[26]) );
  DFFRHQXL array_look_back_reg_3__2_ ( .D(n1538), .CK(clk), .RN(rst_n), .Q(
        array_look_back[38]) );
  DFFRHQXL array_look_back_reg_4__2_ ( .D(n1537), .CK(clk), .RN(rst_n), .Q(
        array_look_back[50]) );
  DFFRHQXL array_look_back_reg_5__2_ ( .D(n1536), .CK(clk), .RN(rst_n), .Q(
        array_look_back[62]) );
  DFFRHQXL array_look_back_reg_6__2_ ( .D(n1535), .CK(clk), .RN(rst_n), .Q(
        array_look_back[74]) );
  DFFRHQXL array_look_back_reg_7__2_ ( .D(n1534), .CK(clk), .RN(rst_n), .Q(
        array_look_back[86]) );
  DFFRHQXL array_look_back_reg_8__2_ ( .D(n1533), .CK(clk), .RN(rst_n), .Q(
        array_look_back[98]) );
  DFFRHQXL array_look_back_reg_9__2_ ( .D(n1532), .CK(clk), .RN(rst_n), .Q(
        array_look_back[110]) );
  DFFRHQXL array_look_back_reg_10__2_ ( .D(n1531), .CK(clk), .RN(rst_n), .Q(
        array_look_back[122]) );
  DFFRHQXL array_look_back_reg_11__2_ ( .D(n1530), .CK(clk), .RN(rst_n), .Q(
        array_look_back[134]) );
  DFFRHQXL array_look_back_reg_11__11_ ( .D(n1681), .CK(clk), .RN(rst_n), .Q(
        array_look_back[143]) );
  DFFRHQXL array_look_back_reg_0__11_ ( .D(n1597), .CK(clk), .RN(rst_n), .Q(
        array_look_back[11]) );
  DFFRHQXL array_look_back_reg_1__11_ ( .D(n1593), .CK(clk), .RN(rst_n), .Q(
        array_look_back[23]) );
  DFFRHQXL array_look_back_reg_2__11_ ( .D(n1589), .CK(clk), .RN(rst_n), .Q(
        array_look_back[35]) );
  DFFRHQXL array_look_back_reg_3__11_ ( .D(n1585), .CK(clk), .RN(rst_n), .Q(
        array_look_back[47]) );
  DFFRHQXL array_look_back_reg_4__11_ ( .D(n1581), .CK(clk), .RN(rst_n), .Q(
        array_look_back[59]) );
  DFFRHQXL array_look_back_reg_5__11_ ( .D(n1577), .CK(clk), .RN(rst_n), .Q(
        array_look_back[71]) );
  DFFRHQXL array_look_back_reg_6__11_ ( .D(n1573), .CK(clk), .RN(rst_n), .Q(
        array_look_back[83]) );
  DFFRHQXL array_look_back_reg_7__11_ ( .D(n1569), .CK(clk), .RN(rst_n), .Q(
        array_look_back[95]) );
  DFFRHQXL array_look_back_reg_8__11_ ( .D(n1565), .CK(clk), .RN(rst_n), .Q(
        array_look_back[107]) );
  DFFRHQXL array_look_back_reg_9__11_ ( .D(n1561), .CK(clk), .RN(rst_n), .Q(
        array_look_back[119]) );
  DFFRHQXL array_look_back_reg_10__11_ ( .D(n1557), .CK(clk), .RN(rst_n), .Q(
        array_look_back[131]) );
  DFFRHQXL array_look_back_reg_0__3_ ( .D(n1553), .CK(clk), .RN(rst_n), .Q(
        array_look_back[3]) );
  DFFRHQXL array_look_back_reg_1__3_ ( .D(n1552), .CK(clk), .RN(rst_n), .Q(
        array_look_back[15]) );
  DFFRHQXL array_look_back_reg_2__3_ ( .D(n1551), .CK(clk), .RN(rst_n), .Q(
        array_look_back[27]) );
  DFFRHQXL array_look_back_reg_3__3_ ( .D(n1550), .CK(clk), .RN(rst_n), .Q(
        array_look_back[39]) );
  DFFRHQXL array_look_back_reg_4__3_ ( .D(n1549), .CK(clk), .RN(rst_n), .Q(
        array_look_back[51]) );
  DFFRHQXL array_look_back_reg_5__3_ ( .D(n1548), .CK(clk), .RN(rst_n), .Q(
        array_look_back[63]) );
  DFFRHQXL array_look_back_reg_6__3_ ( .D(n1547), .CK(clk), .RN(rst_n), .Q(
        array_look_back[75]) );
  DFFRHQXL array_look_back_reg_7__3_ ( .D(n1546), .CK(clk), .RN(rst_n), .Q(
        array_look_back[87]) );
  DFFRHQXL array_look_back_reg_8__3_ ( .D(n1545), .CK(clk), .RN(rst_n), .Q(
        array_look_back[99]) );
  DFFRHQXL array_look_back_reg_9__3_ ( .D(n1544), .CK(clk), .RN(rst_n), .Q(
        array_look_back[111]) );
  DFFRHQXL array_look_back_reg_10__3_ ( .D(n1543), .CK(clk), .RN(rst_n), .Q(
        array_look_back[123]) );
  DFFRHQXL array_look_back_reg_11__3_ ( .D(n1542), .CK(clk), .RN(rst_n), .Q(
        array_look_back[135]) );
  DFFRHQXL array_look_back_reg_0__6_ ( .D(n1493), .CK(clk), .RN(rst_n), .Q(
        array_look_back[6]) );
  DFFRHQXL array_look_back_reg_1__6_ ( .D(n1492), .CK(clk), .RN(rst_n), .Q(
        array_look_back[18]) );
  DFFRHQXL array_look_back_reg_2__6_ ( .D(n1491), .CK(clk), .RN(rst_n), .Q(
        array_look_back[30]) );
  DFFRHQXL array_look_back_reg_3__6_ ( .D(n1490), .CK(clk), .RN(rst_n), .Q(
        array_look_back[42]) );
  DFFRHQXL array_look_back_reg_4__6_ ( .D(n1489), .CK(clk), .RN(rst_n), .Q(
        array_look_back[54]) );
  DFFRHQXL array_look_back_reg_5__6_ ( .D(n1488), .CK(clk), .RN(rst_n), .Q(
        array_look_back[66]) );
  DFFRHQXL array_look_back_reg_6__6_ ( .D(n1487), .CK(clk), .RN(rst_n), .Q(
        array_look_back[78]) );
  DFFRHQXL array_look_back_reg_7__6_ ( .D(n1486), .CK(clk), .RN(rst_n), .Q(
        array_look_back[90]) );
  DFFRHQXL array_look_back_reg_8__6_ ( .D(n1485), .CK(clk), .RN(rst_n), .Q(
        array_look_back[102]) );
  DFFRHQXL array_look_back_reg_9__6_ ( .D(n1484), .CK(clk), .RN(rst_n), .Q(
        array_look_back[114]) );
  DFFRHQXL array_look_back_reg_10__6_ ( .D(n1483), .CK(clk), .RN(rst_n), .Q(
        array_look_back[126]) );
  DFFRHQXL array_look_back_reg_11__6_ ( .D(n1482), .CK(clk), .RN(rst_n), .Q(
        array_look_back[138]) );
  DFFRHQXL array_look_back_reg_0__0_ ( .D(n1517), .CK(clk), .RN(rst_n), .Q(
        array_look_back[0]) );
  DFFRHQXL array_look_back_reg_1__0_ ( .D(n1516), .CK(clk), .RN(rst_n), .Q(
        array_look_back[12]) );
  DFFRHQXL array_look_back_reg_2__0_ ( .D(n1515), .CK(clk), .RN(rst_n), .Q(
        array_look_back[24]) );
  DFFRHQXL array_look_back_reg_3__0_ ( .D(n1514), .CK(clk), .RN(rst_n), .Q(
        array_look_back[36]) );
  DFFRHQXL array_look_back_reg_4__0_ ( .D(n1513), .CK(clk), .RN(rst_n), .Q(
        array_look_back[48]) );
  DFFRHQXL array_look_back_reg_5__0_ ( .D(n1512), .CK(clk), .RN(rst_n), .Q(
        array_look_back[60]) );
  DFFRHQXL array_look_back_reg_6__0_ ( .D(n1511), .CK(clk), .RN(rst_n), .Q(
        array_look_back[72]) );
  DFFRHQXL array_look_back_reg_7__0_ ( .D(n1510), .CK(clk), .RN(rst_n), .Q(
        array_look_back[84]) );
  DFFRHQXL array_look_back_reg_8__0_ ( .D(n1509), .CK(clk), .RN(rst_n), .Q(
        array_look_back[96]) );
  DFFRHQXL array_look_back_reg_9__0_ ( .D(n1508), .CK(clk), .RN(rst_n), .Q(
        array_look_back[108]) );
  DFFRHQXL array_look_back_reg_10__0_ ( .D(n1507), .CK(clk), .RN(rst_n), .Q(
        array_look_back[120]) );
  DFFRHQXL array_look_back_reg_11__0_ ( .D(n1506), .CK(clk), .RN(rst_n), .Q(
        array_look_back[132]) );
  DFFRHQXL array_look_back_reg_0__1_ ( .D(n1529), .CK(clk), .RN(rst_n), .Q(
        array_look_back[1]) );
  DFFRHQXL array_look_back_reg_1__1_ ( .D(n1528), .CK(clk), .RN(rst_n), .Q(
        array_look_back[13]) );
  DFFRHQXL array_look_back_reg_2__1_ ( .D(n1527), .CK(clk), .RN(rst_n), .Q(
        array_look_back[25]) );
  DFFRHQXL array_look_back_reg_3__1_ ( .D(n1526), .CK(clk), .RN(rst_n), .Q(
        array_look_back[37]) );
  DFFRHQXL array_look_back_reg_4__1_ ( .D(n1525), .CK(clk), .RN(rst_n), .Q(
        array_look_back[49]) );
  DFFRHQXL array_look_back_reg_5__1_ ( .D(n1524), .CK(clk), .RN(rst_n), .Q(
        array_look_back[61]) );
  DFFRHQXL array_look_back_reg_6__1_ ( .D(n1523), .CK(clk), .RN(rst_n), .Q(
        array_look_back[73]) );
  DFFRHQXL array_look_back_reg_7__1_ ( .D(n1522), .CK(clk), .RN(rst_n), .Q(
        array_look_back[85]) );
  DFFRHQXL array_look_back_reg_8__1_ ( .D(n1521), .CK(clk), .RN(rst_n), .Q(
        array_look_back[97]) );
  DFFRHQXL array_look_back_reg_9__1_ ( .D(n1520), .CK(clk), .RN(rst_n), .Q(
        array_look_back[109]) );
  DFFRHQXL array_look_back_reg_10__1_ ( .D(n1519), .CK(clk), .RN(rst_n), .Q(
        array_look_back[121]) );
  DFFRHQXL array_look_back_reg_11__1_ ( .D(n1518), .CK(clk), .RN(rst_n), .Q(
        array_look_back[133]) );
  DFFRHQXL array_look_back_reg_0__5_ ( .D(n1481), .CK(clk), .RN(rst_n), .Q(
        array_look_back[5]) );
  DFFRHQXL array_look_back_reg_1__5_ ( .D(n1480), .CK(clk), .RN(rst_n), .Q(
        array_look_back[17]) );
  DFFRHQXL array_look_back_reg_2__5_ ( .D(n1479), .CK(clk), .RN(rst_n), .Q(
        array_look_back[29]) );
  DFFRHQXL array_look_back_reg_3__5_ ( .D(n1478), .CK(clk), .RN(rst_n), .Q(
        array_look_back[41]) );
  DFFRHQXL array_look_back_reg_4__5_ ( .D(n1477), .CK(clk), .RN(rst_n), .Q(
        array_look_back[53]) );
  DFFRHQXL array_look_back_reg_5__5_ ( .D(n1476), .CK(clk), .RN(rst_n), .Q(
        array_look_back[65]) );
  DFFRHQXL array_look_back_reg_6__5_ ( .D(n1475), .CK(clk), .RN(rst_n), .Q(
        array_look_back[77]) );
  DFFRHQXL array_look_back_reg_7__5_ ( .D(n1474), .CK(clk), .RN(rst_n), .Q(
        array_look_back[89]) );
  DFFRHQXL array_look_back_reg_8__5_ ( .D(n1473), .CK(clk), .RN(rst_n), .Q(
        array_look_back[101]) );
  DFFRHQXL array_look_back_reg_9__5_ ( .D(n1472), .CK(clk), .RN(rst_n), .Q(
        array_look_back[113]) );
  DFFRHQXL array_look_back_reg_10__5_ ( .D(n1471), .CK(clk), .RN(rst_n), .Q(
        array_look_back[125]) );
  DFFRHQXL array_look_back_reg_11__5_ ( .D(n1470), .CK(clk), .RN(rst_n), .Q(
        array_look_back[137]) );
  DFFRHQXL y_array_reg_1_ ( .D(n1405), .CK(clk), .RN(rst_n), .Q(y_array[1]) );
  DFFRHQXL y_array_reg_11_ ( .D(n1457), .CK(clk), .RN(rst_n), .Q(y_array[11])
         );
  DFFRHQXL y_array_reg_9_ ( .D(n1455), .CK(clk), .RN(rst_n), .Q(y_array[9]) );
  DFFRHQXL y_array_reg_10_ ( .D(n1456), .CK(clk), .RN(rst_n), .Q(y_array[10])
         );
  DFFRHQXL y_array_reg_8_ ( .D(n1454), .CK(clk), .RN(rst_n), .Q(y_array[8]) );
  DFFRHQXL y_array_reg_3_ ( .D(n1407), .CK(clk), .RN(rst_n), .Q(y_array[3]) );
  DFFRHQXL y_array_reg_2_ ( .D(n1406), .CK(clk), .RN(rst_n), .Q(y_array[2]) );
  DFFRHQXL y_array_reg_6_ ( .D(n1402), .CK(clk), .RN(rst_n), .Q(y_array[6]) );
  DFFRHQXL count_out_reg_3_ ( .D(N6085), .CK(clk), .RN(rst_n), .Q(count_out[3]) );
  DFFHQX1 row_store_reg_0__0_ ( .D(n1395), .CK(clk), .Q(row_store[0]) );
  DFFHQX1 row_store_reg_0__1_ ( .D(n1394), .CK(clk), .Q(row_store[1]) );
  DFFHQX1 row_store_reg_0__2_ ( .D(n1393), .CK(clk), .Q(row_store[2]) );
  DFFHQX1 row_store_reg_0__3_ ( .D(n1392), .CK(clk), .Q(row_store[3]) );
  DFFSX1 out_valid_reg ( .D(n3086), .CK(clk), .SN(rst_n), .QN(out_valid) );
  DFFSX1 count_reg_2_ ( .D(n1661), .CK(clk), .SN(rst_n), .QN(n3084) );
  DFFSX1 count_reg_0_ ( .D(n1663), .CK(clk), .SN(rst_n), .QN(n3083) );
  DFFSX1 count_reg_3_ ( .D(n1662), .CK(clk), .SN(rst_n), .Q(count[3]) );
  DFFSX1 count_reg_1_ ( .D(n1660), .CK(clk), .SN(rst_n), .Q(count[1]) );
  DFFRX1 count_out_reg_0_ ( .D(N6082), .CK(clk), .RN(rst_n), .Q(count_out[0]), 
        .QN(n3085) );
  DFFRHQXL out_reg_3_ ( .D(n1399), .CK(clk), .RN(rst_n), .Q(out[3]) );
  DFFRHQXL out_reg_2_ ( .D(n1398), .CK(clk), .RN(rst_n), .Q(out[2]) );
  DFFRHQXL out_reg_1_ ( .D(n1397), .CK(clk), .RN(rst_n), .Q(out[1]) );
  DFFRHQXL out_reg_0_ ( .D(n1396), .CK(clk), .RN(rst_n), .Q(out[0]) );
  DFFRHQX1 x_reg_3_ ( .D(n1680), .CK(clk), .RN(rst_n), .Q(N4586) );
  DFFRHQX1 x_reg_2_ ( .D(n1615), .CK(clk), .RN(rst_n), .Q(x[2]) );
  NOR2X1 U1686 ( .A(count_out[0]), .B(n3086), .Y(N6082) );
  NOR2X1 U1687 ( .A(n3044), .B(n3043), .Y(n3074) );
  NOR2X1 U1688 ( .A(n2484), .B(n2768), .Y(n2623) );
  NOR2X1 U1689 ( .A(n2797), .B(n2732), .Y(n2739) );
  NOR2X1 U1690 ( .A(n2796), .B(n2795), .Y(n2816) );
  NOR2X1 U1691 ( .A(array_in[7]), .B(n2078), .Y(n2080) );
  AND4X2 U1692 ( .A(n3036), .B(n3035), .C(n3034), .D(n3033), .Y(n3037) );
  AND4X2 U1693 ( .A(n3018), .B(n3017), .C(n3016), .D(n3015), .Y(n3019) );
  AND4X2 U1694 ( .A(n3002), .B(n3001), .C(n3000), .D(n2999), .Y(n3003) );
  AND4X2 U1695 ( .A(n3066), .B(n3065), .C(n3064), .D(n3063), .Y(n3068) );
  NOR2X1 U1696 ( .A(row[0]), .B(n2550), .Y(n2380) );
  NOR2X1 U1697 ( .A(n2517), .B(n2692), .Y(n2185) );
  AOI32X1 U1698 ( .A0(n2438), .A1(n2574), .A2(n2577), .B0(n2760), .B1(n2574), 
        .Y(n2499) );
  NOR2X1 U1699 ( .A(n2788), .B(n2789), .Y(n2774) );
  NOR2X1 U1700 ( .A(n3007), .B(n2661), .Y(n2377) );
  NOR2X1 U1701 ( .A(n2059), .B(n2058), .Y(n2047) );
  NOR2X1 U1702 ( .A(n2222), .B(n2534), .Y(n2531) );
  NOR2X1 U1703 ( .A(n2105), .B(n2034), .Y(n2052) );
  NOR2X1 U1704 ( .A(n2452), .B(n2451), .Y(n2664) );
  NOR2X1 U1705 ( .A(n2458), .B(n2454), .Y(n2675) );
  NOR2X1 U1706 ( .A(current_state[1]), .B(n2024), .Y(n2046) );
  NOR2X1 U1707 ( .A(n2717), .B(n2685), .Y(n2493) );
  NOR2X1 U1708 ( .A(n2346), .B(n2345), .Y(n2350) );
  NOR2X1 U1709 ( .A(n2024), .B(n2023), .Y(n2528) );
  NOR2X1 U1710 ( .A(count_out[2]), .B(n2829), .Y(n3058) );
  NOR2X1 U1711 ( .A(count_out[2]), .B(n2834), .Y(n3053) );
  AND4X2 U1712 ( .A(n2337), .B(n2321), .C(n2320), .D(n2319), .Y(n2322) );
  NOR2X1 U1713 ( .A(n2827), .B(n2831), .Y(n3052) );
  NOR2X1 U1714 ( .A(count_out[3]), .B(n1692), .Y(n3059) );
  AND4X2 U1715 ( .A(n2318), .B(n2317), .C(n2316), .D(n2315), .Y(n2319) );
  NOR2X1 U1716 ( .A(n2128), .B(n2133), .Y(n2123) );
  NOR2X1 U1717 ( .A(count_out[1]), .B(count_out[3]), .Y(n2830) );
  NOR2X1 U1718 ( .A(n2139), .B(n2144), .Y(n2147) );
  AND4X2 U1719 ( .A(n2278), .B(n2277), .C(n2276), .D(n2275), .Y(n2279) );
  AND4X2 U1720 ( .A(n1937), .B(n1936), .C(n1935), .D(n1934), .Y(n2144) );
  NOR2X1 U1721 ( .A(n1771), .B(n1956), .Y(n1792) );
  NOR2X1 U1722 ( .A(n1938), .B(n1989), .Y(n1955) );
  NOR2X1 U1723 ( .A(n1836), .B(n1861), .Y(n1837) );
  NOR2X1 U1724 ( .A(add_array[13]), .B(array_look_back[46]), .Y(n1859) );
  NOR2X1 U1725 ( .A(n1960), .B(n1959), .Y(n1965) );
  NOR2X1 U1726 ( .A(array_look_back[1]), .B(add_array[1]), .Y(n1892) );
  NOR2X1 U1727 ( .A(n2207), .B(n2197), .Y(n2310) );
  NOR2X1 U1728 ( .A(n2212), .B(n2220), .Y(n2313) );
  NOR2X1 U1729 ( .A(n1911), .B(n2632), .Y(n1957) );
  NOR2X1 U1730 ( .A(n2464), .B(n1864), .Y(n1968) );
  NOR2X1 U1731 ( .A(n2304), .B(n2309), .Y(n2101) );
  NOR2X1 U1732 ( .A(x[1]), .B(n2027), .Y(n2029) );
  NOR2X1 U1733 ( .A(n2098), .B(n2017), .Y(n2056) );
  NAND2X1 U1734 ( .A(n2464), .B(n1972), .Y(n2563) );
  INVX2 U1735 ( .A(n1846), .Y(n1958) );
  INVX2 U1736 ( .A(n1951), .Y(n2011) );
  NAND2X1 U1737 ( .A(n2207), .B(n2441), .Y(n2220) );
  INVXL U1738 ( .A(n1911), .Y(n2116) );
  INVXL U1739 ( .A(n2572), .Y(n2423) );
  AOI222XL U1740 ( .A0(n2818), .A1(n2708), .B0(n2707), .B1(n2817), .C0(n2814), 
        .C1(n2706), .Y(n2709) );
  INVX2 U1741 ( .A(n2499), .Y(n2576) );
  NAND3X1 U1742 ( .A(n2329), .B(n2343), .C(n2325), .Y(n2349) );
  OR2XL U1743 ( .A(n2339), .B(n2345), .Y(n2335) );
  INVX2 U1744 ( .A(n2570), .Y(n2178) );
  INVX1 U1745 ( .A(n2398), .Y(n2562) );
  INVX1 U1746 ( .A(n2379), .Y(n2557) );
  INVX2 U1747 ( .A(n2760), .Y(n2425) );
  INVX2 U1748 ( .A(n2692), .Y(n2699) );
  INVX1 U1749 ( .A(n2472), .Y(n2679) );
  INVX1 U1750 ( .A(n2463), .Y(n2683) );
  NOR2BX1 U1751 ( .AN(n2014), .B(n2013), .Y(n2309) );
  INVXL U1752 ( .A(n2096), .Y(n2010) );
  NAND2X1 U1753 ( .A(n1931), .B(n1958), .Y(n2575) );
  OR2X1 U1754 ( .A(array_in[1]), .B(n2029), .Y(n2095) );
  INVX1 U1755 ( .A(n1908), .Y(n1964) );
  NAND2X1 U1756 ( .A(n2685), .B(x[2]), .Y(n1846) );
  INVX2 U1757 ( .A(x[1]), .Y(n2471) );
  INVX2 U1758 ( .A(N4586), .Y(n2685) );
  INVX2 U1759 ( .A(in_valid), .Y(n2168) );
  MXI2XL U1760 ( .A(n2822), .B(n2722), .S0(n2721), .Y(n1425) );
  MXI2XL U1761 ( .A(n2822), .B(n2751), .S0(n2750), .Y(n1417) );
  MXI2XL U1762 ( .A(n2822), .B(n2758), .S0(n2757), .Y(n1415) );
  MXI2XL U1763 ( .A(n2822), .B(n2710), .S0(n2709), .Y(n1427) );
  MXI2XL U1764 ( .A(n2822), .B(n2749), .S0(n2748), .Y(n1418) );
  MXI2XL U1765 ( .A(n2822), .B(n2729), .S0(n2728), .Y(n1423) );
  MXI2XL U1766 ( .A(n2822), .B(n2694), .S0(n2693), .Y(n1429) );
  MXI2XL U1767 ( .A(n2822), .B(n2808), .S0(n2807), .Y(n1410) );
  NOR2X1 U1768 ( .A(n2744), .B(n2655), .Y(n2510) );
  NOR2X1 U1769 ( .A(n2744), .B(n2647), .Y(n2476) );
  OAI21XL U1770 ( .A0(n2582), .A1(n2581), .B0(n2792), .Y(n2599) );
  OAI31XL U1771 ( .A0(n2744), .A1(n2518), .A2(n2760), .B0(n2792), .Y(n2630) );
  AND2XL U1772 ( .A(n2696), .B(n2783), .Y(n2811) );
  OAI2BB1X1 U1773 ( .A0N(n2793), .A1N(n2759), .B0(n2792), .Y(n2708) );
  OAI21XL U1774 ( .A0(n2604), .A1(n2581), .B0(n2792), .Y(n2635) );
  OAI21XL U1775 ( .A0(n2760), .A1(n2490), .B0(n2792), .Y(n2613) );
  OAI2BB1X1 U1776 ( .A0N(n2794), .A1N(n2793), .B0(n2792), .Y(n2819) );
  OAI21XL U1777 ( .A0(n2760), .A1(n2656), .B0(n2792), .Y(n2640) );
  OAI2BB1XL U1778 ( .A0N(n2695), .A1N(n2703), .B0(n2792), .Y(n2775) );
  OAI31XL U1779 ( .A0(n2440), .A1(n2670), .A2(n2659), .B0(n2591), .Y(n2507) );
  NOR2X1 U1780 ( .A(n2413), .B(n2412), .Y(n2415) );
  AOI2BB1XL U1781 ( .A0N(n2452), .A1N(n2453), .B0(n2451), .Y(n2603) );
  NOR2X1 U1782 ( .A(n2390), .B(n2416), .Y(n2392) );
  NOR2X1 U1783 ( .A(n2377), .B(n2376), .Y(n2378) );
  NOR2X1 U1784 ( .A(n2403), .B(n2416), .Y(n2405) );
  OAI2BB1XL U1785 ( .A0N(n2703), .A1N(n2702), .B0(n2792), .Y(n2771) );
  NOR2X1 U1786 ( .A(n2357), .B(n2356), .Y(n2359) );
  NOR2X1 U1787 ( .A(n2397), .B(n2416), .Y(n2399) );
  NOR2X1 U1788 ( .A(n2417), .B(n2416), .Y(n2418) );
  OAI2BB1XL U1789 ( .A0N(n2445), .A1N(n2660), .B0(n2670), .Y(n2591) );
  NOR2X1 U1790 ( .A(n2397), .B(n2410), .Y(n2367) );
  AOI2BB1XL U1791 ( .A0N(n2449), .A1N(n2450), .B0(n2448), .Y(n2453) );
  NOR2X1 U1792 ( .A(n2403), .B(n2410), .Y(n2383) );
  NOR2X1 U1793 ( .A(n2377), .B(n2360), .Y(n2352) );
  NOR2BXL U1794 ( .AN(n2444), .B(n2443), .Y(n2670) );
  NOR2X1 U1795 ( .A(n2662), .B(n2439), .Y(n2443) );
  NAND2XL U1796 ( .A(n2439), .B(n2662), .Y(n2444) );
  NOR2X1 U1797 ( .A(n2660), .B(n2659), .Y(n2671) );
  NOR2X1 U1798 ( .A(n3007), .B(n2439), .Y(n2371) );
  NOR2X1 U1799 ( .A(n2441), .B(n2666), .Y(n2452) );
  AOI211X1 U1800 ( .A0(n2343), .A1(n2342), .B0(n2341), .C0(n2340), .Y(n2659)
         );
  NOR2X1 U1801 ( .A(n2340), .B(n2330), .Y(n2439) );
  NOR2X1 U1802 ( .A(n2449), .B(n2448), .Y(n2669) );
  NOR2X1 U1803 ( .A(n2447), .B(n2667), .Y(n2451) );
  NOR2X1 U1804 ( .A(n2663), .B(n2446), .Y(n2448) );
  OAI211XL U1805 ( .A0(n2327), .A1(n2349), .B0(n2326), .C0(n2325), .Y(n2340)
         );
  NOR2X1 U1806 ( .A(n2349), .B(n2344), .Y(n2447) );
  NOR2X1 U1807 ( .A(n2207), .B(n2442), .Y(n2449) );
  NAND2BXL U1808 ( .AN(n2335), .B(n2338), .Y(n2323) );
  OAI21X1 U1809 ( .A0(n2517), .A1(n2760), .B0(n2576), .Y(n2515) );
  NOR2X1 U1810 ( .A(n2349), .B(n2346), .Y(n2338) );
  OAI2BB1XL U1811 ( .A0N(n2329), .A1N(n2328), .B0(n2343), .Y(n2330) );
  OAI2BB1X1 U1812 ( .A0N(n2426), .A1N(n2425), .B0(n2574), .Y(n2436) );
  AND2X2 U1813 ( .A(n2334), .B(n2332), .Y(n2329) );
  NAND3XL U1814 ( .A(n2274), .B(n2273), .C(n2272), .Y(n2339) );
  AOI211X1 U1815 ( .A0(array_look_back[22]), .A1(n2313), .B0(n2253), .C0(n2252), .Y(n2343) );
  NOR2X1 U1816 ( .A(n2765), .B(n2778), .Y(n2782) );
  NAND3XL U1817 ( .A(n2281), .B(n2280), .C(n2279), .Y(n2345) );
  AOI21X1 U1818 ( .A0(n2179), .A1(n2425), .B0(n2178), .Y(n2572) );
  NAND4XL U1819 ( .A(n2251), .B(n2250), .C(n2249), .D(n2248), .Y(n2252) );
  OAI2BB1XL U1820 ( .A0N(array_look_back[19]), .A1N(n2313), .B0(n2226), .Y(
        n2232) );
  NAND4XL U1821 ( .A(n2230), .B(n2229), .C(n2228), .D(n2227), .Y(n2231) );
  OAI2BB1XL U1822 ( .A0N(array_look_back[106]), .A1N(n2312), .B0(n2247), .Y(
        n2253) );
  OAI2BB1XL U1823 ( .A0N(array_look_back[133]), .A1N(n2304), .B0(n2296), .Y(
        n2302) );
  OAI2BB1XL U1824 ( .A0N(array_look_back[23]), .A1N(n2313), .B0(n2254), .Y(
        n2260) );
  NAND4XL U1825 ( .A(n2258), .B(n2257), .C(n2256), .D(n2255), .Y(n2259) );
  NAND4XL U1826 ( .A(n2286), .B(n2285), .C(n2284), .D(n2283), .Y(n2287) );
  NOR2X1 U1827 ( .A(n2718), .B(n2747), .Y(n2725) );
  OAI2BB1XL U1828 ( .A0N(array_look_back[102]), .A1N(n2312), .B0(n2282), .Y(
        n2288) );
  NOR2X1 U1829 ( .A(n2797), .B(n2747), .Y(n2754) );
  OAI2BB1XL U1830 ( .A0N(array_look_back[98]), .A1N(n2312), .B0(n2289), .Y(
        n2295) );
  NOR2X1 U1831 ( .A(n2765), .B(n2705), .Y(n2809) );
  NOR2X1 U1832 ( .A(n2763), .B(n2762), .Y(n2798) );
  NOR2X1 U1833 ( .A(n2610), .B(n2479), .Y(n2645) );
  NOR2X1 U1834 ( .A(n2692), .B(n2777), .Y(n2804) );
  INVX1 U1835 ( .A(n2351), .Y(n2556) );
  INVX1 U1836 ( .A(n2419), .Y(n2579) );
  INVX1 U1837 ( .A(n2357), .Y(n2564) );
  NOR2X1 U1838 ( .A(n2583), .B(n2494), .Y(n2633) );
  INVX1 U1839 ( .A(n2362), .Y(n2555) );
  NOR2X1 U1840 ( .A(n2610), .B(n2583), .Y(n2597) );
  NOR2X1 U1841 ( .A(n2718), .B(n2732), .Y(n2706) );
  INVX1 U1842 ( .A(n2372), .Y(n2554) );
  AOI21X1 U1843 ( .A0(n2425), .A1(n2167), .B0(n2166), .Y(n2570) );
  INVX1 U1844 ( .A(n2391), .Y(n2567) );
  AOI2BB1XL U1845 ( .A0N(x[1]), .A1N(n2156), .B0(n2160), .Y(n2561) );
  NOR2X1 U1846 ( .A(n2686), .B(n2593), .Y(n2611) );
  NOR2X1 U1847 ( .A(n2145), .B(n2150), .Y(n2351) );
  NOR2X1 U1848 ( .A(n2145), .B(n2152), .Y(n2357) );
  NOR2X1 U1849 ( .A(n2594), .B(n2593), .Y(n2653) );
  INVX1 U1850 ( .A(n2565), .Y(n2166) );
  NAND2XL U1851 ( .A(n2660), .B(n2662), .Y(n2197) );
  NOR2X1 U1852 ( .A(n2161), .B(n2159), .Y(n2398) );
  AOI2BB1XL U1853 ( .A0N(n2171), .A1N(n2692), .B0(n2552), .Y(n2173) );
  NOR2X1 U1854 ( .A(n2202), .B(n2692), .Y(n2204) );
  NOR2X1 U1855 ( .A(n2566), .B(n2692), .Y(n2213) );
  NOR2X1 U1856 ( .A(n2563), .B(n2692), .Y(n2217) );
  NOR2X1 U1857 ( .A(n2463), .B(n2154), .Y(n2413) );
  NOR2X1 U1858 ( .A(n2692), .B(n2797), .Y(n2764) );
  NOR2X1 U1859 ( .A(n2580), .B(n2692), .Y(n2189) );
  NOR2X1 U1860 ( .A(n2571), .B(n2692), .Y(n2175) );
  NOR2X1 U1861 ( .A(n2683), .B(n2154), .Y(n2366) );
  NOR2X1 U1862 ( .A(n2573), .B(n2692), .Y(n2182) );
  OAI211X1 U1863 ( .A0(n2022), .A1(n2021), .B0(n2054), .C0(n2020), .Y(n2662)
         );
  NOR2X1 U1864 ( .A(n2575), .B(n2692), .Y(n2209) );
  NOR2X1 U1865 ( .A(n2438), .B(n2692), .Y(n2194) );
  NOR2X1 U1866 ( .A(n2158), .B(n2148), .Y(n2404) );
  NOR2X1 U1867 ( .A(n2577), .B(n2692), .Y(n2199) );
  AOI2BB1XL U1868 ( .A0N(n2081), .A1N(n2016), .B0(n2015), .Y(n2054) );
  NOR2X1 U1869 ( .A(n2153), .B(n2148), .Y(n2384) );
  NOR2X1 U1870 ( .A(n2680), .B(n2679), .Y(n2687) );
  NAND2BX1 U1871 ( .AN(n2025), .B(n2528), .Y(n2692) );
  INVXL U1872 ( .A(n2101), .Y(n2015) );
  NOR2X1 U1873 ( .A(n2463), .B(n2684), .Y(n2025) );
  NOR2X1 U1874 ( .A(n2144), .B(n2143), .Y(n2472) );
  NAND2X1 U1875 ( .A(n1995), .B(n1994), .Y(n2684) );
  NOR2X1 U1876 ( .A(n2469), .B(n2471), .Y(n2462) );
  NOR2X1 U1877 ( .A(n2304), .B(n2081), .Y(n2441) );
  OAI2BB1X1 U1878 ( .A0N(n1995), .A1N(n1993), .B0(n1994), .Y(n2463) );
  NOR2X1 U1879 ( .A(n2125), .B(n2124), .Y(n2469) );
  NOR2X1 U1880 ( .A(n2124), .B(n2146), .Y(n1994) );
  INVX1 U1881 ( .A(n2147), .Y(n2124) );
  NAND2BXL U1882 ( .AN(n2022), .B(n2021), .Y(n2102) );
  NOR2X1 U1883 ( .A(n2121), .B(n2120), .Y(n1995) );
  INVX1 U1884 ( .A(n2055), .Y(n2099) );
  NOR4XL U1885 ( .A(n1834), .B(n1833), .C(n1832), .D(n1831), .Y(n2128) );
  NOR4XL U1886 ( .A(n1855), .B(n1854), .C(n1853), .D(n1852), .Y(n2133) );
  OAI211XL U1887 ( .A0(array_in[7]), .A1(n2685), .B0(n2014), .C0(n2016), .Y(
        n2055) );
  AOI211X1 U1888 ( .A0(n2010), .A1(n2048), .B0(n2307), .C0(n2009), .Y(n2014)
         );
  AND4X2 U1889 ( .A(n1928), .B(n1906), .C(n1905), .D(n1904), .Y(n2139) );
  INVX1 U1890 ( .A(n1986), .Y(n1928) );
  NOR2X1 U1891 ( .A(n2032), .B(n2008), .Y(n2096) );
  NOR2X1 U1892 ( .A(array_in[5]), .B(n2026), .Y(n2098) );
  NOR2X1 U1893 ( .A(n2087), .B(array_in[9]), .Y(n2090) );
  AND4X2 U1894 ( .A(n1872), .B(n1871), .C(n1870), .D(n1869), .Y(n1873) );
  NOR2X1 U1895 ( .A(n2796), .B(n2768), .Y(n2787) );
  NOR2X1 U1896 ( .A(n1836), .B(n1771), .Y(n1752) );
  NOR2X1 U1897 ( .A(n2006), .B(n2078), .Y(n2026) );
  NOR2X1 U1898 ( .A(n1828), .B(n1938), .Y(n1770) );
  OAI2BB1XL U1899 ( .A0N(n2533), .A1N(n2569), .B0(n2095), .Y(n2012) );
  INVXL U1900 ( .A(n2202), .Y(n2008) );
  NOR2X1 U1901 ( .A(array_in[8]), .B(n2563), .Y(n2009) );
  NOR2X1 U1902 ( .A(n2698), .B(n2704), .Y(n2810) );
  NOR2X1 U1903 ( .A(n1863), .B(n1827), .Y(n1830) );
  NOR2X1 U1904 ( .A(n1863), .B(n1835), .Y(n1838) );
  NOR2X1 U1905 ( .A(n2788), .B(n2704), .Y(n2817) );
  AND4X2 U1906 ( .A(n1707), .B(n1706), .C(n1705), .D(n1704), .Y(n1708) );
  NOR2X1 U1907 ( .A(n2396), .B(n2395), .Y(n2406) );
  NOR2X1 U1908 ( .A(n3081), .B(n2549), .Y(n2363) );
  NOR2X1 U1909 ( .A(n1863), .B(n1789), .Y(n1735) );
  NOR2X1 U1910 ( .A(row[3]), .B(n2549), .Y(n2385) );
  NOR2X1 U1911 ( .A(n2491), .B(n2592), .Y(n2612) );
  NOR2X1 U1912 ( .A(n2395), .B(n2551), .Y(n2420) );
  NOR2X1 U1913 ( .A(n2675), .B(n2592), .Y(n2651) );
  NOR2X1 U1914 ( .A(n2586), .B(n2606), .Y(n2598) );
  NOR2X1 U1915 ( .A(n2795), .B(n2731), .Y(n2707) );
  NOR2X1 U1916 ( .A(n2607), .B(n2606), .Y(n2622) );
  NOR2X1 U1917 ( .A(n2746), .B(n2731), .Y(n2740) );
  NAND2X2 U1918 ( .A(n2464), .B(n1967), .Y(n2202) );
  INVX1 U1919 ( .A(n2573), .Y(n2179) );
  NOR2X1 U1920 ( .A(n3007), .B(n3072), .Y(n3076) );
  INVX1 U1921 ( .A(n2571), .Y(n2167) );
  NOR2X1 U1922 ( .A(array_in[1]), .B(n2569), .Y(n2092) );
  INVX1 U1923 ( .A(n2566), .Y(n2149) );
  NOR2X1 U1924 ( .A(n2789), .B(n2698), .Y(n2769) );
  NOR2X1 U1925 ( .A(n2584), .B(n2586), .Y(n2519) );
  NOR2X1 U1926 ( .A(n2464), .B(n1964), .Y(n1973) );
  NOR2X2 U1927 ( .A(n2685), .B(n1864), .Y(n1967) );
  NOR2X1 U1928 ( .A(n2169), .B(n2168), .Y(n2697) );
  NOR2X2 U1929 ( .A(n2685), .B(n2011), .Y(n1969) );
  NOR2X1 U1930 ( .A(n2027), .B(array_in[4]), .Y(n2085) );
  NOR2X1 U1931 ( .A(current_state[2]), .B(n2046), .Y(n2110) );
  NOR2X1 U1932 ( .A(n2168), .B(n3007), .Y(n2532) );
  INVX1 U1933 ( .A(n2007), .Y(n1887) );
  NAND2X1 U1934 ( .A(n2685), .B(n2464), .Y(n2027) );
  NOR2X2 U1935 ( .A(n2680), .B(n2471), .Y(n1951) );
  NOR2X1 U1936 ( .A(n2680), .B(x[1]), .Y(n1908) );
  NOR2X1 U1937 ( .A(n2103), .B(n2985), .Y(n2038) );
  NAND2XL U1938 ( .A(n2065), .B(N4586), .Y(n2013) );
  NOR2X1 U1939 ( .A(n2711), .B(n2222), .Y(n2188) );
  NOR2X1 U1940 ( .A(n2460), .B(n2459), .Y(n2673) );
  INVX2 U1941 ( .A(x[0]), .Y(n2680) );
  NOR2X1 U1942 ( .A(x[0]), .B(x[1]), .Y(n1931) );
  INVX2 U1943 ( .A(x[2]), .Y(n2464) );
  NOR2X1 U1944 ( .A(row[2]), .B(n3079), .Y(n2407) );
  NOR2X1 U1945 ( .A(row[1]), .B(n2456), .Y(n2454) );
  NOR2X1 U1946 ( .A(col[2]), .B(n2672), .Y(n2170) );
  NOR2X1 U1947 ( .A(col[2]), .B(n3080), .Y(n2460) );
  NOR2X1 U1948 ( .A(n3078), .B(col[0]), .Y(n2457) );
  NOR2X1 U1949 ( .A(col[1]), .B(n3079), .Y(n2458) );
  NOR2X1 U1950 ( .A(row[2]), .B(n2455), .Y(n2459) );
  NOR2X1 U1951 ( .A(n2672), .B(n3078), .Y(n2674) );
  INVX1 U1952 ( .A(col[3]), .Y(n2711) );
  NAND2X1 U1953 ( .A(n2018), .B(n1908), .Y(n2566) );
  NAND2X1 U1954 ( .A(n2018), .B(n1951), .Y(n2573) );
  NAND2X1 U1955 ( .A(n2018), .B(n1987), .Y(n2571) );
  INVX2 U1956 ( .A(n2027), .Y(n2018) );
  NAND4BXL U1957 ( .AN(n2323), .B(n2331), .C(n2324), .D(n2322), .Y(n2347) );
  AOI22XL U1958 ( .A0(array_look_back[132]), .A1(n2304), .B0(
        array_look_back[36]), .B1(n2303), .Y(n2321) );
  AOI22XL U1959 ( .A0(array_look_back[48]), .A1(n2306), .B0(
        array_look_back[60]), .B1(n2305), .Y(n2320) );
  AOI2BB1XL U1960 ( .A0N(n2324), .A1N(n2323), .B0(n2344), .Y(n2326) );
  AOI22XL U1961 ( .A0(array_look_back[125]), .A1(n2307), .B0(
        array_look_back[77]), .B1(n2310), .Y(n2274) );
  AOI22XL U1962 ( .A0(array_look_back[101]), .A1(n2312), .B0(
        array_look_back[113]), .B1(n2308), .Y(n2273) );
  AOI22XL U1963 ( .A0(array_look_back[59]), .A1(n2306), .B0(
        array_look_back[143]), .B1(n2304), .Y(n2254) );
  AOI211XL U1964 ( .A0(array_look_back[139]), .A1(n2304), .B0(n2232), .C0(
        n2231), .Y(n2327) );
  AOI22XL U1965 ( .A0(array_look_back[7]), .A1(n2314), .B0(array_look_back[55]), .B1(n2306), .Y(n2226) );
  AOI32XL U1966 ( .A0(n1819), .A1(n1818), .A2(n1848), .B0(n2011), .B1(n1818), 
        .Y(n1834) );
  NAND4XL U1967 ( .A(n1823), .B(n1822), .C(n1821), .D(n1820), .Y(n1833) );
  OAI211XL U1968 ( .A0(n1826), .A1(n2902), .B0(n1825), .C0(n1824), .Y(n1832)
         );
  OAI211XL U1969 ( .A0(n1735), .A1(n2011), .B0(n1734), .C0(n1733), .Y(n2129)
         );
  OAI21XL U1970 ( .A0(n1827), .A1(n1828), .B0(n1908), .Y(n1733) );
  NOR4XL U1971 ( .A(n1986), .B(n1728), .C(n1727), .D(n1726), .Y(n1734) );
  OAI22XL U1972 ( .A0(n1838), .A1(n1964), .B0(n1837), .B1(n2117), .Y(n1855) );
  NAND4XL U1973 ( .A(n1842), .B(n1841), .C(n1840), .D(n1839), .Y(n1854) );
  OAI211XL U1974 ( .A0(n2569), .A1(n2151), .B0(n1844), .C0(n1843), .Y(n1853)
         );
  OAI211XL U1975 ( .A0(n2680), .A1(n1880), .B0(n1928), .C0(n1879), .Y(n2131)
         );
  OAI32XL U1976 ( .A0(x[1]), .A1(n1862), .A2(n1861), .B0(n1860), .B1(n2471), 
        .Y(n1880) );
  AOI211XL U1977 ( .A0(n2149), .A1(array_look_back[22]), .B0(n1878), .C0(n1877), .Y(n1879) );
  OAI211XL U1978 ( .A0(n1859), .A1(n2027), .B0(n1858), .C0(n1857), .Y(n1860)
         );
  AOI22XL U1979 ( .A0(array_look_back[80]), .A1(n2310), .B0(
        array_look_back[128]), .B1(n2307), .Y(n2246) );
  AOI211XL U1980 ( .A0(array_look_back[6]), .A1(n2314), .B0(n2288), .C0(n2287), 
        .Y(n2333) );
  AOI22XL U1981 ( .A0(array_look_back[42]), .A1(n2303), .B0(
        array_look_back[126]), .B1(n2307), .Y(n2285) );
  AOI211XL U1982 ( .A0(array_look_back[14]), .A1(n2313), .B0(n2295), .C0(n2294), .Y(n2331) );
  NAND4XL U1983 ( .A(n2293), .B(n2292), .C(n2291), .D(n2290), .Y(n2294) );
  AOI22XL U1984 ( .A0(array_look_back[134]), .A1(n2304), .B0(
        array_look_back[122]), .B1(n2307), .Y(n2292) );
  AOI22XL U1985 ( .A0(array_look_back[81]), .A1(n2310), .B0(
        array_look_back[129]), .B1(n2307), .Y(n2239) );
  AOI211XL U1986 ( .A0(array_look_back[13]), .A1(n2313), .B0(n2302), .C0(n2301), .Y(n2337) );
  NAND4XL U1987 ( .A(n2300), .B(n2299), .C(n2298), .D(n2297), .Y(n2301) );
  AOI22XL U1988 ( .A0(array_look_back[1]), .A1(n2314), .B0(array_look_back[49]), .B1(n2306), .Y(n2296) );
  AOI22XL U1989 ( .A0(array_look_back[10]), .A1(n2314), .B0(
        array_look_back[70]), .B1(n2305), .Y(n2247) );
  OAI211XL U1990 ( .A0(n2018), .A1(array_in[3]), .B0(n2056), .C0(n2099), .Y(
        n2022) );
  NAND2XL U1991 ( .A(n2985), .B(n2086), .Y(n2021) );
  AOI21XL U1992 ( .A0(n2438), .A1(n2026), .B0(array_in[4]), .Y(n2017) );
  NAND2XL U1993 ( .A(x[2]), .B(n1951), .Y(n2005) );
  NAND2XL U1994 ( .A(n2007), .B(n2171), .Y(n2032) );
  NAND2XL U1995 ( .A(n2685), .B(n2005), .Y(n2078) );
  NAND2XL U1996 ( .A(array_in[9]), .B(array_in[8]), .Y(n2048) );
  INVXL U1997 ( .A(n1952), .Y(n1772) );
  NAND2XL U1998 ( .A(n1795), .B(n1794), .Y(n1835) );
  AOI22XL U1999 ( .A0(n2018), .A1(sub_array[3]), .B0(n1958), .B1(sub_array[7]), 
        .Y(n1795) );
  AOI22XL U2000 ( .A0(n1887), .A1(sub_array[15]), .B0(n2116), .B1(
        sub_array[11]), .Y(n1794) );
  AOI22XL U2001 ( .A0(n1973), .A1(array_look_back[61]), .B0(add_array[9]), 
        .B1(n1970), .Y(n1899) );
  NAND2XL U2002 ( .A(x[2]), .B(n1931), .Y(n1826) );
  NAND2XL U2003 ( .A(n1886), .B(n1885), .Y(n1959) );
  AOI22XL U2004 ( .A0(n2018), .A1(add_array[3]), .B0(n1958), .B1(add_array[7]), 
        .Y(n1886) );
  AOI22XL U2005 ( .A0(n1887), .A1(add_array[15]), .B0(n2116), .B1(
        add_array[11]), .Y(n1885) );
  INVXL U2006 ( .A(n1918), .Y(n1971) );
  AOI2BB1XL U2007 ( .A0N(array_look_back[11]), .A1N(sub_array[0]), .B0(n2569), 
        .Y(n1802) );
  INVXL U2008 ( .A(n1835), .Y(n1867) );
  INVXL U2009 ( .A(n1826), .Y(n1966) );
  AOI211XL U2010 ( .A0(n1931), .A1(n1988), .B0(n1930), .C0(n1929), .Y(n1935)
         );
  OAI211XL U2011 ( .A0(n1912), .A1(n1911), .B0(n1910), .C0(n1909), .Y(n1930)
         );
  NAND4XL U2012 ( .A(n1928), .B(n1927), .C(n1926), .D(n1925), .Y(n1929) );
  OAI211XL U2013 ( .A0(n1752), .A1(n2011), .B0(n1751), .C0(n1750), .Y(n2127)
         );
  OAI2BB1XL U2014 ( .A0N(n1819), .A1N(n1775), .B0(n1908), .Y(n1750) );
  NOR4XL U2015 ( .A(n1986), .B(n1749), .C(n1748), .D(n1747), .Y(n1751) );
  OAI211XL U2016 ( .A0(n1792), .A1(n1964), .B0(n1791), .C0(n1790), .Y(n2134)
         );
  OAI21XL U2017 ( .A0(n1789), .A1(n1989), .B0(n1931), .Y(n1790) );
  NOR4XL U2018 ( .A(n1986), .B(n1786), .C(n1785), .D(n1784), .Y(n1791) );
  AOI22XL U2019 ( .A0(array_look_back[124]), .A1(n2307), .B0(
        array_look_back[76]), .B1(n2310), .Y(n2281) );
  AOI22XL U2020 ( .A0(array_look_back[100]), .A1(n2312), .B0(
        array_look_back[112]), .B1(n2308), .Y(n2280) );
  NAND2XL U2021 ( .A(n2339), .B(n2338), .Y(n2348) );
  OAI32XL U2022 ( .A0(n2679), .A1(n2462), .A2(x[0]), .B0(x[1]), .B1(n2470), 
        .Y(n2467) );
  NAND2XL U2023 ( .A(x[1]), .B(n2469), .Y(n2681) );
  INVXL U2024 ( .A(n2659), .Y(n2445) );
  NAND2XL U2025 ( .A(n2137), .B(n2134), .Y(n2120) );
  NAND2XL U2026 ( .A(n2126), .B(n2141), .Y(n2146) );
  NAND2XL U2027 ( .A(n2129), .B(n2127), .Y(n2121) );
  OAI211XL U2028 ( .A0(n1992), .A1(n2011), .B0(n1991), .C0(n1990), .Y(n2141)
         );
  AOI211XL U2029 ( .A0(sub_array[16]), .A1(n1958), .B0(n1957), .C0(n1956), .Y(
        n1992) );
  OAI21XL U2030 ( .A0(n1989), .A1(n1988), .B0(n1987), .Y(n1990) );
  NOR4XL U2031 ( .A(n1986), .B(n1985), .C(n1984), .D(n1983), .Y(n1991) );
  AOI22XL U2032 ( .A0(n1969), .A1(array_look_back[132]), .B0(n1966), .B1(
        array_look_back[48]), .Y(n1936) );
  OAI2BB1XL U2033 ( .A0N(n1933), .A1N(n1932), .B0(x[2]), .Y(n1934) );
  AOI22XL U2034 ( .A0(n1968), .A1(array_look_back[72]), .B0(n2424), .B1(
        add_array[4]), .Y(n1937) );
  AOI22XL U2035 ( .A0(sub_array[16]), .A1(n2006), .B0(n2426), .B1(add_array[6]), .Y(n1906) );
  AOI22XL U2036 ( .A0(n1951), .A1(n1884), .B0(n1931), .B1(n1960), .Y(n1905) );
  NOR4XL U2037 ( .A(n1903), .B(n1902), .C(n1901), .D(n1900), .Y(n1904) );
  INVXL U2038 ( .A(n2129), .Y(n2130) );
  OAI211XL U2039 ( .A0(n1770), .A1(n2011), .B0(n1769), .C0(n1768), .Y(n2137)
         );
  OAI21XL U2040 ( .A0(n1789), .A1(n1952), .B0(n1908), .Y(n1768) );
  NOR4XL U2041 ( .A(n1986), .B(n1767), .C(n1766), .D(n1765), .Y(n1769) );
  OAI211XL U2042 ( .A0(n1955), .A1(n1964), .B0(n1954), .C0(n1953), .Y(n2126)
         );
  OAI21XL U2043 ( .A0(n1952), .A1(n1988), .B0(n1951), .Y(n1953) );
  NOR4XL U2044 ( .A(n1986), .B(n1950), .C(n1949), .D(n1948), .Y(n1954) );
  NAND2XL U2045 ( .A(n2528), .B(n2472), .Y(n2153) );
  INVXL U2046 ( .A(n2469), .Y(n2470) );
  INVXL U2047 ( .A(n2569), .Y(n2119) );
  NAND2XL U2048 ( .A(n2469), .B(n2472), .Y(n2145) );
  INVXL U2049 ( .A(n2575), .Y(n2424) );
  NAND2XL U2050 ( .A(n2659), .B(n2792), .Y(n2355) );
  AOI222XL U2051 ( .A0(row[1]), .A1(col[1]), .B0(row[1]), .B1(n2674), .C0(
        col[1]), .C1(n2674), .Y(n2676) );
  INVXL U2052 ( .A(n2702), .Y(n2695) );
  OAI2BB1XL U2053 ( .A0N(n2682), .A1N(n2687), .B0(n2681), .Y(n2689) );
  NAND2XL U2054 ( .A(n2767), .B(n2766), .Y(n2796) );
  MXI2XL U2055 ( .A(x[0]), .B(n2680), .S0(n2472), .Y(n2797) );
  XOR2XL U2056 ( .A(n2713), .B(n2712), .Y(n2766) );
  NAND2XL U2057 ( .A(n2763), .B(n2762), .Y(n2747) );
  XOR2XL U2058 ( .A(n2671), .B(n2670), .Y(n2702) );
  XNOR2XL U2059 ( .A(n2669), .B(n2668), .Y(n2703) );
  INVXL U2060 ( .A(n2788), .Y(n2698) );
  NAND2XL U2061 ( .A(n2697), .B(n2789), .Y(n2704) );
  AND2XL U2062 ( .A(n2745), .B(n2744), .Y(n2793) );
  NAND2XL U2063 ( .A(n2713), .B(n2678), .Y(n2731) );
  NOR2X1 U2064 ( .A(col[3]), .B(row[3]), .Y(n2678) );
  XOR2XL U2065 ( .A(n2483), .B(n2712), .Y(n2584) );
  NOR3XL U2066 ( .A(n2603), .B(n2760), .C(n2489), .Y(n2480) );
  NAND2XL U2067 ( .A(n2583), .B(n2609), .Y(n2479) );
  OAI2BB1XL U2068 ( .A0N(n2483), .A1N(n2482), .B0(n2481), .Y(n2585) );
  INVXL U2069 ( .A(n2582), .Y(n2604) );
  AOI21XL U2070 ( .A0(n2468), .A1(n2492), .B0(n2493), .Y(n2609) );
  INVXL U2071 ( .A(n2586), .Y(n2607) );
  XOR2XL U2072 ( .A(n2660), .B(n2445), .Y(n2744) );
  AOI22XL U2073 ( .A0(n2472), .A1(n2594), .B0(n2686), .B1(n2679), .Y(n2475) );
  XOR2XL U2074 ( .A(n2664), .B(n2453), .Y(n2582) );
  NAND2XL U2075 ( .A(n2603), .B(n2489), .Y(n2581) );
  XOR2XL U2076 ( .A(n2673), .B(n2461), .Y(n2586) );
  NAND2XL U2077 ( .A(n2585), .B(n2584), .Y(n2606) );
  XOR2XL U2078 ( .A(n2714), .B(n2492), .Y(n2610) );
  NOR2X2 U2079 ( .A(n2685), .B(n1964), .Y(n1972) );
  AOI21XL U2080 ( .A0(n2097), .A1(n2019), .B0(n2307), .Y(n2020) );
  NOR4XL U2081 ( .A(n2018), .B(n2017), .C(array_in[3]), .D(n2055), .Y(n2097)
         );
  INVXL U2082 ( .A(n2413), .Y(n2568) );
  INVXL U2083 ( .A(n2404), .Y(n2559) );
  AOI21X1 U2084 ( .A0(n2424), .A1(n2425), .B0(n2423), .Y(n2574) );
  AND2XL U2085 ( .A(n2798), .B(n2797), .Y(n2815) );
  XOR2XL U2086 ( .A(n2675), .B(n2674), .Y(n2788) );
  OAI21XL U2087 ( .A0(n2695), .A1(n2703), .B0(n2792), .Y(n2783) );
  INVXL U2088 ( .A(n2770), .Y(n2781) );
  XOR2XL U2089 ( .A(n2673), .B(n2676), .Y(n2789) );
  NAND2XL U2090 ( .A(n2798), .B(n2764), .Y(n2778) );
  NAND2XL U2091 ( .A(n2770), .B(n2765), .Y(n2777) );
  XOR2XL U2092 ( .A(n2689), .B(n2688), .Y(n2770) );
  NOR3XL U2093 ( .A(n2767), .B(n2746), .C(n2766), .Y(n2755) );
  NOR3XL U2094 ( .A(n2767), .B(n2766), .C(n2795), .Y(n2726) );
  OAI31XL U2095 ( .A0(n2703), .A1(n2702), .A2(n2760), .B0(n2792), .Y(n2818) );
  NOR2BXL U2096 ( .AN(n2765), .B(n2705), .Y(n2814) );
  AND2X1 U2097 ( .A(n2771), .B(n2696), .Y(n2801) );
  AND2XL U2098 ( .A(n2697), .B(n2769), .Y(n2800) );
  NOR3XL U2099 ( .A(n2765), .B(n2781), .C(n2692), .Y(n2799) );
  INVXL U2100 ( .A(n2507), .Y(n2518) );
  NOR3XL U2101 ( .A(n2607), .B(n2584), .C(n2585), .Y(n2650) );
  NAND2XL U2102 ( .A(n2744), .B(n2591), .Y(n2656) );
  NAND2XL U2103 ( .A(n2744), .B(n2507), .Y(n2490) );
  NAND2XL U2104 ( .A(n2582), .B(n2480), .Y(n2655) );
  NOR2BXL U2105 ( .AN(n2610), .B(n2479), .Y(n2652) );
  OAI31X1 U2106 ( .A0(n2603), .A1(n2602), .A2(n2604), .B0(n2792), .Y(n2641) );
  NOR2BXL U2107 ( .AN(n2519), .B(n2585), .Y(n2639) );
  AND2XL U2108 ( .A(n2609), .B(n2608), .Y(n2638) );
  AND2XL U2109 ( .A(n2519), .B(n2585), .Y(n2634) );
  NAND2XL U2110 ( .A(n2493), .B(n2492), .Y(n2494) );
  INVXL U2111 ( .A(n2605), .Y(n2625) );
  AOI31XL U2112 ( .A0(n2604), .A1(n2603), .A2(n2602), .B0(n3007), .Y(n2605) );
  NOR3XL U2113 ( .A(n2610), .B(n2609), .C(n2608), .Y(n2621) );
  OAI31XL U2114 ( .A0(n2744), .A1(n2760), .A2(n2507), .B0(n2792), .Y(n2624) );
  NOR2BXL U2115 ( .AN(n2764), .B(n2475), .Y(n2620) );
  NOR2BXL U2116 ( .AN(n2484), .B(n2768), .Y(n2629) );
  AND2XL U2117 ( .A(n2764), .B(n2475), .Y(n2628) );
  NAND2XL U2118 ( .A(n2697), .B(n2531), .Y(n3077) );
  NAND2XL U2119 ( .A(n2685), .B(n1961), .Y(n2517) );
  NAND2XL U2120 ( .A(n1931), .B(n2116), .Y(n2580) );
  NOR3XL U2121 ( .A(n2307), .B(n2096), .C(array_in[9]), .Y(n2308) );
  OAI21XL U2122 ( .A0(n2216), .A1(n2534), .B0(n2792), .Y(n2539) );
  OAI21XL U2123 ( .A0(n2216), .A1(n2181), .B0(n2792), .Y(n2541) );
  OAI31XL U2124 ( .A0(col[1]), .A1(n2711), .A2(n2216), .B0(n2792), .Y(n2547)
         );
  OAI21XL U2125 ( .A0(n2222), .A1(n2198), .B0(n2792), .Y(n2540) );
  OAI21XL U2126 ( .A0(n2198), .A1(n2208), .B0(n2792), .Y(n2544) );
  OAI31XL U2127 ( .A0(n2396), .A1(n2208), .A2(n2534), .B0(n2792), .Y(n2542) );
  OAI31XL U2128 ( .A0(n2396), .A1(n2193), .A2(n2534), .B0(n2792), .Y(n2543) );
  OAI21XL U2129 ( .A0(n2198), .A1(n2193), .B0(n2792), .Y(n2545) );
  OAI21XL U2130 ( .A0(col[1]), .A1(n2203), .B0(n2792), .Y(n2546) );
  OAI21XL U2131 ( .A0(n2456), .A1(n2203), .B0(n2792), .Y(n2548) );
  NAND2X1 U2132 ( .A(n2025), .B(n2528), .Y(n2760) );
  AOI22XL U2133 ( .A0(n2699), .A1(n2037), .B0(n2047), .B1(n2036), .Y(n2114) );
  INVXL U2134 ( .A(col[1]), .Y(n2456) );
  OAI31XL U2135 ( .A0(add_array[3]), .A1(sub_array[14]), .A2(
        array_look_back[36]), .B0(n2179), .Y(n1922) );
  OAI31XL U2136 ( .A0(add_array[2]), .A1(sub_array[13]), .A2(
        array_look_back[24]), .B0(n2167), .Y(n1921) );
  OAI31XL U2137 ( .A0(add_array[1]), .A1(sub_array[12]), .A2(
        array_look_back[12]), .B0(n2149), .Y(n1920) );
  AOI31XL U2138 ( .A0(n1958), .A1(n1951), .A2(sub_array[18]), .B0(n1915), .Y(
        n1917) );
  AOI2BB1XL U2139 ( .A0N(array_look_back[0]), .A1N(add_array[0]), .B0(n2569), 
        .Y(n1915) );
  INVXL U2140 ( .A(n1836), .Y(n1817) );
  INVXL U2141 ( .A(n1827), .Y(n1845) );
  AOI22XL U2142 ( .A0(array_look_back[96]), .A1(n2312), .B0(
        array_look_back[24]), .B1(n2311), .Y(n2316) );
  NAND2XL U2143 ( .A(n1714), .B(n1713), .Y(n1849) );
  AOI22XL U2144 ( .A0(n2018), .A1(sub_array[4]), .B0(n1958), .B1(sub_array[8]), 
        .Y(n1714) );
  AOI22XL U2145 ( .A0(n1887), .A1(sub_array[16]), .B0(n2116), .B1(
        sub_array[12]), .Y(n1713) );
  AOI22XL U2146 ( .A0(array_look_back[89]), .A1(n2309), .B0(
        array_look_back[65]), .B1(n2305), .Y(n2269) );
  AOI22XL U2147 ( .A0(array_look_back[5]), .A1(n2314), .B0(array_look_back[53]), .B1(n2306), .Y(n2271) );
  AOI22XL U2148 ( .A0(array_look_back[29]), .A1(n2311), .B0(
        array_look_back[41]), .B1(n2303), .Y(n2268) );
  AOI22XL U2149 ( .A0(array_look_back[17]), .A1(n2313), .B0(
        array_look_back[137]), .B1(n2304), .Y(n2270) );
  AOI22XL U2150 ( .A0(array_look_back[95]), .A1(n2309), .B0(
        array_look_back[71]), .B1(n2305), .Y(n2256) );
  AOI22XL U2151 ( .A0(array_look_back[107]), .A1(n2312), .B0(
        array_look_back[119]), .B1(n2308), .Y(n2257) );
  AOI22XL U2152 ( .A0(array_look_back[47]), .A1(n2303), .B0(
        array_look_back[35]), .B1(n2311), .Y(n2255) );
  AOI22XL U2153 ( .A0(array_look_back[131]), .A1(n2307), .B0(
        array_look_back[83]), .B1(n2310), .Y(n2258) );
  AOI22XL U2154 ( .A0(array_look_back[103]), .A1(n2312), .B0(
        array_look_back[115]), .B1(n2308), .Y(n2229) );
  AOI22XL U2155 ( .A0(array_look_back[91]), .A1(n2309), .B0(
        array_look_back[67]), .B1(n2305), .Y(n2228) );
  AOI22XL U2156 ( .A0(array_look_back[127]), .A1(n2307), .B0(
        array_look_back[79]), .B1(n2310), .Y(n2230) );
  AOI22XL U2157 ( .A0(array_look_back[31]), .A1(n2311), .B0(
        array_look_back[43]), .B1(n2303), .Y(n2227) );
  AOI22XL U2158 ( .A0(array_look_back[99]), .A1(n2312), .B0(
        array_look_back[111]), .B1(n2308), .Y(n2264) );
  AOI22XL U2159 ( .A0(array_look_back[63]), .A1(n2305), .B0(
        array_look_back[87]), .B1(n2309), .Y(n2263) );
  AOI22XL U2160 ( .A0(array_look_back[27]), .A1(n2311), .B0(
        array_look_back[39]), .B1(n2303), .Y(n2262) );
  AOI22XL U2161 ( .A0(array_look_back[75]), .A1(n2310), .B0(
        array_look_back[123]), .B1(n2307), .Y(n2265) );
  INVXL U2162 ( .A(n1938), .Y(n1982) );
  INVXL U2163 ( .A(n1895), .Y(n1979) );
  AOI22XL U2164 ( .A0(n1971), .A1(array_look_back[98]), .B0(add_array[10]), 
        .B1(n1970), .Y(n1975) );
  AOI211XL U2165 ( .A0(n1961), .A1(array_look_back[84]), .B0(n1924), .C0(n1923), .Y(n1925) );
  OAI211XL U2166 ( .A0(n1919), .A1(n1918), .B0(n1917), .C0(n1916), .Y(n1924)
         );
  NAND3XL U2167 ( .A(n1922), .B(n1921), .C(n1920), .Y(n1923) );
  AOI2BB1XL U2168 ( .A0N(n2720), .A1N(x[2]), .B0(array_look_back[96]), .Y(
        n1919) );
  AOI22XL U2169 ( .A0(add_array[9]), .A1(n2087), .B0(add_array[7]), .B1(n1913), 
        .Y(n1927) );
  INVXL U2170 ( .A(n2517), .Y(n1913) );
  AOI211XL U2171 ( .A0(add_array[10]), .A1(n2008), .B0(y_array[0]), .C0(n1914), 
        .Y(n1926) );
  AOI21XL U2172 ( .A0(n2617), .A1(n2738), .B0(n2438), .Y(n1914) );
  AOI22XL U2173 ( .A0(n1967), .A1(array_look_back[120]), .B0(add_array[11]), 
        .B1(n2157), .Y(n1909) );
  AOI22XL U2174 ( .A0(n1973), .A1(array_look_back[60]), .B0(n1972), .B1(
        array_look_back[108]), .Y(n1910) );
  NAND2XL U2175 ( .A(n1931), .B(n1887), .Y(n1895) );
  AOI21XL U2176 ( .A0(n2119), .A1(array_look_back[8]), .B0(y_array[8]), .Y(
        n1824) );
  AOI22XL U2177 ( .A0(n2149), .A1(array_look_back[20]), .B0(n2167), .B1(
        array_look_back[32]), .Y(n1825) );
  AOI22XL U2178 ( .A0(n2179), .A1(array_look_back[44]), .B0(n1961), .B1(
        array_look_back[92]), .Y(n1821) );
  AOI22XL U2179 ( .A0(n1969), .A1(array_look_back[140]), .B0(n1968), .B1(
        array_look_back[80]), .Y(n1822) );
  OAI2BB1XL U2180 ( .A0N(n1858), .A1N(n1817), .B0(n1908), .Y(n1818) );
  OAI211XL U2181 ( .A0(n1830), .A1(n1864), .B0(n1928), .C0(n1829), .Y(n1831)
         );
  OAI21XL U2182 ( .A0(n1828), .A1(n1835), .B0(n1931), .Y(n1829) );
  OAI211XL U2183 ( .A0(n1817), .A1(n1864), .B0(n1718), .C0(n1717), .Y(n1728)
         );
  OAI2BB1XL U2184 ( .A0N(n1858), .A1N(n1775), .B0(n1931), .Y(n1717) );
  AOI22XL U2185 ( .A0(n2119), .A1(array_look_back[7]), .B0(n1969), .B1(
        array_look_back[139]), .Y(n1718) );
  OAI211XL U2186 ( .A0(n1819), .A1(n1864), .B0(n1725), .C0(n1724), .Y(n1726)
         );
  AOI22XL U2187 ( .A0(n2149), .A1(array_look_back[19]), .B0(n2179), .B1(
        array_look_back[43]), .Y(n1724) );
  NAND4BXL U2188 ( .AN(y_array[7]), .B(n1721), .C(n1720), .D(n1719), .Y(n1727)
         );
  AOI22XL U2189 ( .A0(n2167), .A1(array_look_back[31]), .B0(n1971), .B1(
        array_look_back[103]), .Y(n1721) );
  AOI22XL U2190 ( .A0(n1967), .A1(array_look_back[127]), .B0(n1968), .B1(
        array_look_back[79]), .Y(n1720) );
  NAND2XL U2191 ( .A(n1701), .B(n1700), .Y(n1863) );
  AOI22XL U2192 ( .A0(n2018), .A1(add_array[10]), .B0(n1958), .B1(
        add_array[14]), .Y(n1701) );
  AOI22XL U2193 ( .A0(n1887), .A1(add_array[22]), .B0(n2116), .B1(
        add_array[18]), .Y(n1700) );
  NAND2XL U2194 ( .A(n1730), .B(n1729), .Y(n1827) );
  AOI22XL U2195 ( .A0(n2018), .A1(sub_array[5]), .B0(n1958), .B1(sub_array[9]), 
        .Y(n1730) );
  AOI22XL U2196 ( .A0(n1887), .A1(sub_array[17]), .B0(n2116), .B1(
        sub_array[13]), .Y(n1729) );
  AOI22XL U2197 ( .A0(n2149), .A1(array_look_back[21]), .B0(n2167), .B1(
        array_look_back[33]), .Y(n1844) );
  OAI211XL U2198 ( .A0(n1851), .A1(n2011), .B0(n1928), .C0(n1850), .Y(n1852)
         );
  INVXL U2199 ( .A(n1847), .Y(n1851) );
  OAI21XL U2200 ( .A0(n1849), .A1(n1862), .B0(n1987), .Y(n1850) );
  OAI211XL U2201 ( .A0(n1846), .A1(n2803), .B0(n1865), .C0(n1845), .Y(n1847)
         );
  NAND2XL U2202 ( .A(n1723), .B(n1722), .Y(n1757) );
  AOI22XL U2203 ( .A0(n2018), .A1(sub_array[6]), .B0(n1958), .B1(sub_array[10]), .Y(n1723) );
  AOI22XL U2204 ( .A0(n1887), .A1(sub_array[18]), .B0(n2116), .B1(
        sub_array[14]), .Y(n1722) );
  OAI211XL U2205 ( .A0(n1772), .A1(n2117), .B0(n1746), .C0(n1745), .Y(n1747)
         );
  AOI22XL U2206 ( .A0(n2179), .A1(array_look_back[42]), .B0(n2167), .B1(
        array_look_back[30]), .Y(n1745) );
  OAI211XL U2207 ( .A0(n1845), .A1(n2117), .B0(n1739), .C0(n1738), .Y(n1749)
         );
  OAI21XL U2208 ( .A0(n1828), .A1(n1789), .B0(n1987), .Y(n1738) );
  AOI22XL U2209 ( .A0(n2119), .A1(array_look_back[6]), .B0(n1968), .B1(
        array_look_back[78]), .Y(n1739) );
  NAND4BXL U2210 ( .AN(y_array[6]), .B(n1742), .C(n1741), .D(n1740), .Y(n1748)
         );
  AOI22XL U2211 ( .A0(n1969), .A1(array_look_back[138]), .B0(n1971), .B1(
        array_look_back[102]), .Y(n1742) );
  AOI22XL U2212 ( .A0(n2149), .A1(array_look_back[18]), .B0(n1967), .B1(
        array_look_back[126]), .Y(n1741) );
  AND2XL U2213 ( .A(n1716), .B(n1715), .Y(n1775) );
  AOI22XL U2214 ( .A0(n2018), .A1(add_array[7]), .B0(n1958), .B1(add_array[11]), .Y(n1716) );
  AOI22XL U2215 ( .A0(n1887), .A1(add_array[19]), .B0(n2116), .B1(
        add_array[15]), .Y(n1715) );
  INVXL U2216 ( .A(n1757), .Y(n1819) );
  NAND2XL U2217 ( .A(n1712), .B(n1711), .Y(n1836) );
  AOI22XL U2218 ( .A0(n2018), .A1(add_array[9]), .B0(n1958), .B1(add_array[13]), .Y(n1712) );
  AOI22XL U2219 ( .A0(n1887), .A1(add_array[21]), .B0(n2116), .B1(
        add_array[17]), .Y(n1711) );
  OAI211XL U2220 ( .A0(n1783), .A1(n2011), .B0(n1782), .C0(n1781), .Y(n1784)
         );
  AOI22XL U2221 ( .A0(n1973), .A1(array_look_back[64]), .B0(n1971), .B1(
        array_look_back[100]), .Y(n1781) );
  AOI22XL U2222 ( .A0(n2119), .A1(array_look_back[4]), .B0(n1969), .B1(
        array_look_back[136]), .Y(n1782) );
  NAND4BXL U2223 ( .AN(y_array[4]), .B(n1778), .C(n1777), .D(n1776), .Y(n1785)
         );
  AOI22XL U2224 ( .A0(n1967), .A1(array_look_back[124]), .B0(n1968), .B1(
        array_look_back[76]), .Y(n1776) );
  AOI22XL U2225 ( .A0(n2179), .A1(array_look_back[40]), .B0(n2167), .B1(
        array_look_back[28]), .Y(n1778) );
  OAI211XL U2226 ( .A0(n1775), .A1(n2011), .B0(n1774), .C0(n1773), .Y(n1786)
         );
  OAI2BB1XL U2227 ( .A0N(n1772), .A1N(n1982), .B0(n1987), .Y(n1773) );
  AOI22XL U2228 ( .A0(n2149), .A1(array_look_back[16]), .B0(n1966), .B1(
        array_look_back[52]), .Y(n1774) );
  NAND2XL U2229 ( .A(n1737), .B(n1736), .Y(n1771) );
  AOI22XL U2230 ( .A0(n2018), .A1(sub_array[8]), .B0(n1958), .B1(sub_array[12]), .Y(n1737) );
  AOI22XL U2231 ( .A0(n1887), .A1(sub_array[20]), .B0(n2116), .B1(
        sub_array[16]), .Y(n1736) );
  AOI22XL U2232 ( .A0(n1966), .A1(x_array[4]), .B0(n1968), .B1(x_array[6]), 
        .Y(n1704) );
  AOI22XL U2233 ( .A0(n1961), .A1(x_array[7]), .B0(n1971), .B1(x_array[8]), 
        .Y(n1705) );
  AOI22XL U2234 ( .A0(n1967), .A1(x_array[10]), .B0(n1973), .B1(x_array[5]), 
        .Y(n1706) );
  AOI22XL U2235 ( .A0(n1972), .A1(x_array[9]), .B0(n1969), .B1(x_array[11]), 
        .Y(n1707) );
  INVXL U2236 ( .A(n1771), .Y(n1947) );
  AOI22XL U2237 ( .A0(array_look_back[108]), .A1(n2308), .B0(
        array_look_back[120]), .B1(n2307), .Y(n2318) );
  AOI22XL U2238 ( .A0(array_look_back[0]), .A1(n2314), .B0(array_look_back[12]), .B1(n2313), .Y(n2315) );
  AOI22XL U2239 ( .A0(array_look_back[72]), .A1(n2310), .B0(
        array_look_back[84]), .B1(n2309), .Y(n2317) );
  AOI22XL U2240 ( .A0(array_look_back[64]), .A1(n2305), .B0(
        array_look_back[88]), .B1(n2309), .Y(n2276) );
  AOI22XL U2241 ( .A0(array_look_back[40]), .A1(n2303), .B0(
        array_look_back[28]), .B1(n2311), .Y(n2275) );
  AOI22XL U2242 ( .A0(array_look_back[52]), .A1(n2306), .B0(array_look_back[4]), .B1(n2314), .Y(n2278) );
  AOI22XL U2243 ( .A0(array_look_back[16]), .A1(n2313), .B0(
        array_look_back[136]), .B1(n2304), .Y(n2277) );
  OAI22XL U2244 ( .A0(n1911), .A1(n2791), .B0(n1846), .B1(n2773), .Y(n1856) );
  NAND2XL U2245 ( .A(n1813), .B(n1812), .Y(n1861) );
  AOI22XL U2246 ( .A0(n2018), .A1(sub_array[2]), .B0(n1958), .B1(sub_array[6]), 
        .Y(n1813) );
  AOI22XL U2247 ( .A0(n1887), .A1(sub_array[14]), .B0(n2116), .B1(
        sub_array[10]), .Y(n1812) );
  INVXL U2248 ( .A(n1849), .Y(n1858) );
  NAND4XL U2249 ( .A(n1876), .B(n1875), .C(n1874), .D(n1873), .Y(n1877) );
  AOI32XL U2250 ( .A0(n1867), .A1(n1866), .A2(n1865), .B0(n1864), .B1(n1866), 
        .Y(n1878) );
  AOI22XL U2251 ( .A0(n1931), .A1(n1863), .B0(n2167), .B1(array_look_back[34]), 
        .Y(n1866) );
  INVXL U2252 ( .A(n1848), .Y(n1862) );
  AOI22XL U2253 ( .A0(array_look_back[20]), .A1(n2313), .B0(
        array_look_back[140]), .B1(n2304), .Y(n2242) );
  AOI22XL U2254 ( .A0(array_look_back[66]), .A1(n2305), .B0(
        array_look_back[18]), .B1(n2313), .Y(n2282) );
  AOI22XL U2255 ( .A0(array_look_back[90]), .A1(n2309), .B0(
        array_look_back[54]), .B1(n2306), .Y(n2284) );
  AOI22XL U2256 ( .A0(array_look_back[138]), .A1(n2304), .B0(
        array_look_back[30]), .B1(n2311), .Y(n2283) );
  AOI22XL U2257 ( .A0(array_look_back[78]), .A1(n2310), .B0(
        array_look_back[114]), .B1(n2308), .Y(n2286) );
  AOI22XL U2258 ( .A0(array_look_back[2]), .A1(n2314), .B0(array_look_back[62]), .B1(n2305), .Y(n2289) );
  AOI22XL U2259 ( .A0(array_look_back[86]), .A1(n2309), .B0(
        array_look_back[50]), .B1(n2306), .Y(n2291) );
  AOI22XL U2260 ( .A0(array_look_back[26]), .A1(n2311), .B0(
        array_look_back[38]), .B1(n2303), .Y(n2290) );
  AOI22XL U2261 ( .A0(array_look_back[74]), .A1(n2310), .B0(
        array_look_back[110]), .B1(n2308), .Y(n2293) );
  AOI22XL U2262 ( .A0(array_look_back[109]), .A1(n2308), .B0(
        array_look_back[97]), .B1(n2312), .Y(n2299) );
  AOI22XL U2263 ( .A0(array_look_back[61]), .A1(n2305), .B0(
        array_look_back[85]), .B1(n2309), .Y(n2298) );
  AOI22XL U2264 ( .A0(array_look_back[37]), .A1(n2303), .B0(
        array_look_back[25]), .B1(n2311), .Y(n2297) );
  AOI22XL U2265 ( .A0(array_look_back[73]), .A1(n2310), .B0(
        array_look_back[121]), .B1(n2307), .Y(n2300) );
  AOI211XL U2266 ( .A0(array_look_back[3]), .A1(n2314), .B0(n2267), .C0(n2266), 
        .Y(n2324) );
  OAI2BB1XL U2267 ( .A0N(array_look_back[15]), .A1N(n2313), .B0(n2261), .Y(
        n2267) );
  NAND4XL U2268 ( .A(n2265), .B(n2264), .C(n2263), .D(n2262), .Y(n2266) );
  AOI22XL U2269 ( .A0(array_look_back[51]), .A1(n2306), .B0(
        array_look_back[135]), .B1(n2304), .Y(n2261) );
  AOI22XL U2270 ( .A0(array_look_back[118]), .A1(n2308), .B0(
        array_look_back[82]), .B1(n2310), .Y(n2251) );
  AOI22XL U2271 ( .A0(array_look_back[130]), .A1(n2307), .B0(
        array_look_back[94]), .B1(n2309), .Y(n2250) );
  NAND2XL U2272 ( .A(n2987), .B(n2078), .Y(n2016) );
  INVXL U2273 ( .A(n2347), .Y(n2344) );
  OAI211XL U2274 ( .A0(n1982), .A1(n2117), .B0(n1981), .C0(n1980), .Y(n1983)
         );
  OAI21XL U2275 ( .A0(sub_array[12]), .A1(array_look_back[38]), .B0(n2179), 
        .Y(n1980) );
  AOI211XL U2276 ( .A0(n1979), .A1(add_array[14]), .B0(y_array[2]), .C0(n1978), 
        .Y(n1981) );
  AOI2BB1XL U2277 ( .A0N(add_array[2]), .A1N(array_look_back[2]), .B0(n2569), 
        .Y(n1978) );
  OAI211XL U2278 ( .A0(n1965), .A1(n1964), .B0(n1963), .C0(n1962), .Y(n1985)
         );
  AOI22XL U2279 ( .A0(n2149), .A1(array_look_back[14]), .B0(n1961), .B1(
        array_look_back[86]), .Y(n1963) );
  AOI22XL U2280 ( .A0(n2167), .A1(array_look_back[26]), .B0(n2424), .B1(
        add_array[6]), .Y(n1962) );
  NAND4XL U2281 ( .A(n1977), .B(n1976), .C(n1975), .D(n1974), .Y(n1984) );
  AOI22XL U2282 ( .A0(n1967), .A1(array_look_back[122]), .B0(n1966), .B1(
        array_look_back[50]), .Y(n1977) );
  AOI22XL U2283 ( .A0(n1973), .A1(array_look_back[62]), .B0(n1972), .B1(
        array_look_back[110]), .Y(n1974) );
  AOI22XL U2284 ( .A0(n1969), .A1(array_look_back[134]), .B0(n1968), .B1(
        array_look_back[74]), .Y(n1976) );
  NAND2XL U2285 ( .A(n1756), .B(n1755), .Y(n1956) );
  AOI22XL U2286 ( .A0(n2018), .A1(add_array[5]), .B0(n1958), .B1(add_array[9]), 
        .Y(n1756) );
  AOI22XL U2287 ( .A0(n1887), .A1(add_array[17]), .B0(n2116), .B1(
        add_array[13]), .Y(n1755) );
  AOI22XL U2288 ( .A0(n1967), .A1(add_array[14]), .B0(n1971), .B1(
        add_array[12]), .Y(n1933) );
  AOI22XL U2289 ( .A0(n1972), .A1(add_array[13]), .B0(n1969), .B1(
        add_array[15]), .Y(n1932) );
  OAI211XL U2290 ( .A0(n1892), .A1(n2569), .B0(n1891), .C0(n1890), .Y(n1902)
         );
  OAI21XL U2291 ( .A0(sub_array[13]), .A1(array_look_back[37]), .B0(n2179), 
        .Y(n1890) );
  OAI211XL U2292 ( .A0(n1895), .A1(n2753), .B0(n1894), .C0(n1893), .Y(n1901)
         );
  AOI22XL U2293 ( .A0(n1966), .A1(array_look_back[49]), .B0(n1968), .B1(
        array_look_back[73]), .Y(n1894) );
  OAI21XL U2294 ( .A0(sub_array[12]), .A1(array_look_back[25]), .B0(n2167), 
        .Y(n1893) );
  NAND4XL U2295 ( .A(n1899), .B(n1898), .C(n1897), .D(n1896), .Y(n1900) );
  AOI22XL U2296 ( .A0(n1961), .A1(array_look_back[85]), .B0(n2424), .B1(
        add_array[5]), .Y(n1897) );
  AOI32XL U2297 ( .A0(n1907), .A1(n1889), .A2(n1888), .B0(n1964), .B1(n1889), 
        .Y(n1903) );
  OAI21XL U2298 ( .A0(n1959), .A1(n1957), .B0(n1987), .Y(n1889) );
  NAND2XL U2299 ( .A(n1780), .B(n1779), .Y(n1960) );
  AOI22XL U2300 ( .A0(n2018), .A1(sub_array[10]), .B0(n1958), .B1(
        sub_array[14]), .Y(n1780) );
  AOI22XL U2301 ( .A0(n1887), .A1(sub_array[22]), .B0(n2116), .B1(
        sub_array[18]), .Y(n1779) );
  NAND2BXL U2302 ( .AN(n1989), .B(n1883), .Y(n1884) );
  AOI22XL U2303 ( .A0(n2116), .A1(sub_array[21]), .B0(n1958), .B1(
        sub_array[17]), .Y(n1883) );
  INVXL U2304 ( .A(n2577), .Y(n2006) );
  OAI211XL U2305 ( .A0(n1947), .A1(n1864), .B0(n1764), .C0(n1763), .Y(n1765)
         );
  AOI22XL U2306 ( .A0(n1968), .A1(array_look_back[77]), .B0(n1961), .B1(
        array_look_back[89]), .Y(n1764) );
  AOI22XL U2307 ( .A0(n2149), .A1(array_look_back[17]), .B0(n2179), .B1(
        array_look_back[41]), .Y(n1763) );
  OAI211XL U2308 ( .A0(n1775), .A1(n1864), .B0(n1759), .C0(n1758), .Y(n1767)
         );
  OAI21XL U2309 ( .A0(n1757), .A1(n1956), .B0(n1931), .Y(n1758) );
  AOI22XL U2310 ( .A0(n2119), .A1(array_look_back[5]), .B0(n1967), .B1(
        array_look_back[125]), .Y(n1759) );
  NAND4BXL U2311 ( .AN(y_array[5]), .B(n1762), .C(n1761), .D(n1760), .Y(n1766)
         );
  AOI22XL U2312 ( .A0(n1972), .A1(array_look_back[113]), .B0(n1966), .B1(
        array_look_back[53]), .Y(n1761) );
  AOI22XL U2313 ( .A0(n1973), .A1(array_look_back[65]), .B0(n1969), .B1(
        array_look_back[137]), .Y(n1760) );
  AOI22XL U2314 ( .A0(n2167), .A1(array_look_back[29]), .B0(n1971), .B1(
        array_look_back[101]), .Y(n1762) );
  NAND2XL U2315 ( .A(n1703), .B(n1702), .Y(n1789) );
  AOI22XL U2316 ( .A0(n2018), .A1(sub_array[7]), .B0(n1958), .B1(sub_array[11]), .Y(n1703) );
  AOI22XL U2317 ( .A0(n1887), .A1(sub_array[19]), .B0(n2116), .B1(
        sub_array[15]), .Y(n1702) );
  NAND2XL U2318 ( .A(n1732), .B(n1731), .Y(n1828) );
  AOI22XL U2319 ( .A0(n2018), .A1(add_array[8]), .B0(n1958), .B1(add_array[12]), .Y(n1732) );
  AOI22XL U2320 ( .A0(n1887), .A1(add_array[20]), .B0(n2116), .B1(
        add_array[16]), .Y(n1731) );
  NAND3X1 U2321 ( .A(n1710), .B(n1709), .C(n1708), .Y(n1986) );
  AOI22XL U2322 ( .A0(n2149), .A1(x_array[1]), .B0(n2179), .B1(x_array[3]), 
        .Y(n1710) );
  AOI22XL U2323 ( .A0(n2119), .A1(x_array[0]), .B0(n2167), .B1(x_array[2]), 
        .Y(n1709) );
  NAND4BXL U2324 ( .AN(y_array[3]), .B(n1944), .C(n1943), .D(n1942), .Y(n1949)
         );
  AOI22XL U2325 ( .A0(n2167), .A1(array_look_back[27]), .B0(n1971), .B1(
        array_look_back[99]), .Y(n1944) );
  AOI22XL U2326 ( .A0(n2179), .A1(array_look_back[39]), .B0(n1966), .B1(
        array_look_back[51]), .Y(n1942) );
  OAI211XL U2327 ( .A0(n1941), .A1(n2117), .B0(n1940), .C0(n1939), .Y(n1950)
         );
  INVXL U2328 ( .A(n1959), .Y(n1941) );
  OAI21XL U2329 ( .A0(n1956), .A1(n1960), .B0(n1987), .Y(n1939) );
  AOI22XL U2330 ( .A0(n2119), .A1(array_look_back[3]), .B0(n1973), .B1(
        array_look_back[63]), .Y(n1940) );
  OAI211XL U2331 ( .A0(n1947), .A1(n2117), .B0(n1946), .C0(n1945), .Y(n1948)
         );
  AOI22XL U2332 ( .A0(n1968), .A1(array_look_back[75]), .B0(n1961), .B1(
        array_look_back[87]), .Y(n1946) );
  AOI22XL U2333 ( .A0(n2149), .A1(array_look_back[15]), .B0(n1972), .B1(
        array_look_back[111]), .Y(n1945) );
  NAND2XL U2334 ( .A(n1744), .B(n1743), .Y(n1952) );
  AOI22XL U2335 ( .A0(n2018), .A1(add_array[6]), .B0(n1958), .B1(add_array[10]), .Y(n1744) );
  AOI22XL U2336 ( .A0(n1887), .A1(add_array[18]), .B0(n2116), .B1(
        add_array[14]), .Y(n1743) );
  INVXL U2337 ( .A(n1907), .Y(n1988) );
  NAND2XL U2338 ( .A(n1754), .B(n1753), .Y(n1938) );
  AOI22XL U2339 ( .A0(n2018), .A1(sub_array[9]), .B0(n1958), .B1(sub_array[13]), .Y(n1754) );
  AOI22XL U2340 ( .A0(n1887), .A1(sub_array[21]), .B0(n2116), .B1(
        sub_array[17]), .Y(n1753) );
  NAND2XL U2341 ( .A(n1788), .B(n1787), .Y(n1989) );
  AOI22XL U2342 ( .A0(n2018), .A1(add_array[4]), .B0(n1958), .B1(add_array[8]), 
        .Y(n1788) );
  AOI22XL U2343 ( .A0(n1887), .A1(add_array[16]), .B0(n2116), .B1(
        add_array[12]), .Y(n1787) );
  NAND2XL U2344 ( .A(n2327), .B(n2333), .Y(n2346) );
  AOI22XL U2345 ( .A0(sub_array[5]), .A1(n2426), .B0(sub_array[8]), .B1(n1970), 
        .Y(n1815) );
  OAI21XL U2346 ( .A0(n1861), .A1(n1856), .B0(n1987), .Y(n1814) );
  AOI22XL U2347 ( .A0(n1961), .A1(array_look_back[95]), .B0(n1971), .B1(
        array_look_back[107]), .Y(n1816) );
  NOR4BXL U2348 ( .AN(n1809), .B(y_array[11]), .C(n1808), .D(n1807), .Y(n1810)
         );
  OAI211XL U2349 ( .A0(n2724), .A1(n2566), .B0(n1800), .C0(n1799), .Y(n1808)
         );
  NAND4XL U2350 ( .A(n1806), .B(n1805), .C(n1804), .D(n1803), .Y(n1807) );
  AOI22XL U2351 ( .A0(n1908), .A1(n1798), .B0(n1951), .B1(n1797), .Y(n1811) );
  INVXL U2352 ( .A(n2447), .Y(n2666) );
  AOI222XL U2353 ( .A0(n2677), .A1(col[2]), .B0(n2677), .B1(row[2]), .C0(
        col[2]), .C1(row[2]), .Y(n2713) );
  INVXL U2354 ( .A(n2676), .Y(n2677) );
  NAND2XL U2355 ( .A(n2482), .B(n2481), .Y(n2712) );
  NAND2XL U2356 ( .A(col[3]), .B(n3081), .Y(n2481) );
  AOI31XL U2357 ( .A0(n2660), .A1(n2445), .A2(n2444), .B0(n2443), .Y(n2450) );
  NAND2XL U2358 ( .A(n2685), .B(n2717), .Y(n2468) );
  NAND2XL U2359 ( .A(n2471), .B(n2470), .Y(n2682) );
  INVXL U2360 ( .A(n2602), .Y(n2489) );
  OAI22XL U2361 ( .A0(n2458), .A1(n2457), .B0(row[1]), .B1(n2456), .Y(n2461)
         );
  NOR2BXL U2362 ( .AN(n2468), .B(n2493), .Y(n2714) );
  INVXL U2363 ( .A(n2014), .Y(n2081) );
  NAND2XL U2364 ( .A(N4586), .B(x[2]), .Y(n2007) );
  NAND2XL U2365 ( .A(n2464), .B(N4586), .Y(n1911) );
  NOR2X1 U2366 ( .A(n2835), .B(n2829), .Y(n3061) );
  NOR2X1 U2367 ( .A(n2526), .B(n2833), .Y(n3056) );
  NOR2X1 U2368 ( .A(count_out[1]), .B(n2831), .Y(n3055) );
  NAND2XL U2369 ( .A(n2679), .B(n2528), .Y(n2158) );
  NAND2XL U2370 ( .A(n2147), .B(n2146), .Y(n2148) );
  OAI31XL U2371 ( .A0(n2447), .A1(n2442), .A2(n2760), .B0(n2792), .Y(n2370) );
  NAND2XL U2372 ( .A(n2717), .B(n2699), .Y(n2150) );
  INVXL U2373 ( .A(n1931), .Y(n2117) );
  OAI21XL U2374 ( .A0(n2331), .A1(n2335), .B0(n2333), .Y(n2328) );
  OAI211XL U2375 ( .A0(n2350), .A1(n2349), .B0(n2348), .C0(n2347), .Y(n2442)
         );
  NAND2XL U2376 ( .A(n2684), .B(n2470), .Y(n2159) );
  OR2XL U2377 ( .A(n2158), .B(n2683), .Y(n2161) );
  NAND2XL U2378 ( .A(n2116), .B(n2696), .Y(n2156) );
  OAI211XL U2379 ( .A0(n1882), .A1(n1881), .B0(n2123), .C0(n2131), .Y(n1993)
         );
  OAI211XL U2380 ( .A0(n1848), .A1(n2117), .B0(n1811), .C0(n1810), .Y(n1882)
         );
  NAND4XL U2381 ( .A(n1928), .B(n1816), .C(n1815), .D(n1814), .Y(n1881) );
  OR2XL U2382 ( .A(n2153), .B(n2159), .Y(n2154) );
  NAND2XL U2383 ( .A(n2466), .B(n2465), .Y(n2688) );
  NAND2XL U2384 ( .A(n2464), .B(n2463), .Y(n2466) );
  NAND2XL U2385 ( .A(x[2]), .B(n2683), .Y(n2465) );
  NAND2XL U2386 ( .A(n2699), .B(n2781), .Y(n2705) );
  NAND2XL U2387 ( .A(n2792), .B(n2760), .Y(n2696) );
  INVXL U2388 ( .A(n2746), .Y(n2795) );
  NAND3XL U2389 ( .A(n2685), .B(n2684), .C(n2715), .Y(n2732) );
  XOR2XL U2390 ( .A(n2687), .B(n2686), .Y(n2765) );
  OAI31XL U2391 ( .A0(n2337), .A1(n2336), .A2(n2335), .B0(n2334), .Y(n2342) );
  NAND3XL U2392 ( .A(n2333), .B(n2332), .C(n2331), .Y(n2336) );
  AOI2BB1XL U2393 ( .A0N(n2459), .A1N(n2461), .B0(n2460), .Y(n2483) );
  NAND2XL U2394 ( .A(row[3]), .B(n2711), .Y(n2482) );
  AOI21XL U2395 ( .A0(n3078), .A1(col[0]), .B0(n2457), .Y(n2746) );
  XOR2XL U2396 ( .A(n2688), .B(n2467), .Y(n2608) );
  NAND2XL U2397 ( .A(n2681), .B(n2682), .Y(n2594) );
  OAI2BB2XL U2398 ( .B0(n2491), .B1(n2457), .A0N(n2457), .A1N(n2491), .Y(n2484) );
  NAND2XL U2399 ( .A(n2697), .B(n2795), .Y(n2768) );
  INVXL U2400 ( .A(n2608), .Y(n2583) );
  INVXL U2401 ( .A(n2675), .Y(n2491) );
  INVXL U2402 ( .A(n2594), .Y(n2686) );
  NAND2XL U2403 ( .A(n2699), .B(n2797), .Y(n2593) );
  NAND2XL U2404 ( .A(n2697), .B(n2170), .Y(n2216) );
  NAND2XL U2405 ( .A(n2697), .B(n2174), .Y(n2198) );
  NAND2XL U2406 ( .A(n2697), .B(n2188), .Y(n2203) );
  NAND2XL U2407 ( .A(n2046), .B(n1998), .Y(n2169) );
  AND2XL U2408 ( .A(n2987), .B(n2026), .Y(n2042) );
  INVXL U2409 ( .A(n2439), .Y(n2661) );
  INVXL U2410 ( .A(n2442), .Y(n2663) );
  NAND2XL U2411 ( .A(n2792), .B(n2445), .Y(n2388) );
  OAI2BB1XL U2412 ( .A0N(n2425), .A1N(n2447), .B0(n2792), .Y(n2389) );
  NAND2XL U2413 ( .A(n3078), .B(n3081), .Y(n2395) );
  INVXL U2414 ( .A(n2120), .Y(n2122) );
  AOI221XL U2415 ( .A0(n2142), .A1(n2141), .B0(n2140), .B1(n2141), .C0(n2139), 
        .Y(n2143) );
  NAND2XL U2416 ( .A(n2683), .B(n2699), .Y(n2152) );
  INVXL U2417 ( .A(col[2]), .Y(n2455) );
  INVXL U2418 ( .A(col[0]), .Y(n2672) );
  INVXL U2419 ( .A(n2181), .Y(n2174) );
  AOI2BB1XL U2420 ( .A0N(n2168), .A1N(n2068), .B0(n3007), .Y(n2067) );
  INVXL U2421 ( .A(n2580), .Y(n1970) );
  NAND2XL U2422 ( .A(N4586), .B(n1931), .Y(n1918) );
  OAI2BB1XL U2423 ( .A0N(array_in[7]), .A1N(n1697), .B0(n2517), .Y(n1699) );
  NOR2X1 U2424 ( .A(n2835), .B(n2834), .Y(n3051) );
  INVXL U2425 ( .A(row[3]), .Y(n3081) );
  INVXL U2426 ( .A(row[2]), .Y(n3080) );
  INVXL U2427 ( .A(row[0]), .Y(n3078) );
  NOR2BXL U2428 ( .AN(rst_n), .B(n3077), .Y(n3082) );
  NOR3XL U2429 ( .A(n2472), .B(n2470), .C(n2152), .Y(n2391) );
  AOI2BB1XL U2430 ( .A0N(n2442), .A1N(n2439), .B0(n3007), .Y(n2403) );
  NOR3XL U2431 ( .A(n2469), .B(n2472), .C(n2150), .Y(n2372) );
  NAND2XL U2432 ( .A(n2370), .B(n2388), .Y(n2376) );
  NOR3XL U2433 ( .A(n2684), .B(n2470), .C(n2161), .Y(n2379) );
  NOR3XL U2434 ( .A(n2469), .B(n2679), .C(n2150), .Y(n2362) );
  NAND2XL U2435 ( .A(n2355), .B(n2370), .Y(n2360) );
  INVXL U2436 ( .A(n2384), .Y(n2558) );
  OAI31XL U2437 ( .A0(n2119), .A1(n2118), .A2(n2760), .B0(n2792), .Y(n2160) );
  AOI2BB1XL U2438 ( .A0N(n2117), .A1N(x[2]), .B0(n2685), .Y(n2118) );
  AOI21XL U2439 ( .A0(n2149), .A1(n2425), .B0(n3007), .Y(n2565) );
  AOI2BB1XL U2440 ( .A0N(n2439), .A1N(n2663), .B0(n3007), .Y(n2390) );
  AOI2BB1XL U2441 ( .A0N(n2661), .A1N(n2442), .B0(n3007), .Y(n2397) );
  NOR2X1 U2442 ( .A(row[1]), .B(row[2]), .Y(n2400) );
  NAND2XL U2443 ( .A(n2578), .B(n2156), .Y(n2164) );
  OAI21XL U2444 ( .A0(n2157), .A1(n2156), .B0(n2561), .Y(n2162) );
  INVXL U2445 ( .A(n2561), .Y(n2155) );
  INVXL U2446 ( .A(n2160), .Y(n2578) );
  NAND2XL U2447 ( .A(n2389), .B(n2355), .Y(n2410) );
  NAND2XL U2448 ( .A(row[2]), .B(n2385), .Y(n2411) );
  AND2X1 U2449 ( .A(n2696), .B(n2775), .Y(n2806) );
  AND2XL U2450 ( .A(n2697), .B(n2774), .Y(n2805) );
  NAND2XL U2451 ( .A(n2480), .B(n2604), .Y(n2647) );
  NOR3XL U2452 ( .A(n2483), .B(n2607), .C(n2482), .Y(n2644) );
  NAND2XL U2453 ( .A(n2484), .B(n2650), .Y(n2485) );
  NAND2XL U2454 ( .A(n2697), .B(n2746), .Y(n2592) );
  NAND2XL U2455 ( .A(n2697), .B(row[2]), .Y(n2551) );
  NAND2XL U2456 ( .A(n2697), .B(row[0]), .Y(n2549) );
  NAND2XL U2457 ( .A(n2697), .B(row[3]), .Y(n2550) );
  OAI31XL U2458 ( .A0(n2456), .A1(n2711), .A2(n2216), .B0(n2792), .Y(n2552) );
  NAND2XL U2459 ( .A(n2697), .B(row[1]), .Y(n2553) );
  NAND2XL U2460 ( .A(n1998), .B(current_state[1]), .Y(n2023) );
  NOR2X1 U2461 ( .A(n2104), .B(n2990), .Y(n2039) );
  NOR2X1 U2462 ( .A(n2043), .B(n2092), .Y(n2045) );
  NOR2X1 U2463 ( .A(n2042), .B(n2028), .Y(n2057) );
  NOR2X1 U2464 ( .A(n2092), .B(n2040), .Y(n2063) );
  NAND2XL U2465 ( .A(n2018), .B(n2011), .Y(n2086) );
  OAI2BB1XL U2466 ( .A0N(n2027), .A1N(n2575), .B0(n2104), .Y(n2084) );
  AOI211XL U2467 ( .A0(n2099), .A1(n2098), .B0(n2097), .C0(n2308), .Y(n2100)
         );
  OAI2BB1XL U2468 ( .A0N(n2107), .A1N(array_in[9]), .B0(array_in[8]), .Y(n2108) );
  AOI2BB1XL U2469 ( .A0N(n2661), .A1N(n2663), .B0(n3007), .Y(n2417) );
  NAND2XL U2470 ( .A(n2389), .B(n2388), .Y(n2416) );
  NOR3XL U2471 ( .A(n2469), .B(n2472), .C(n2152), .Y(n2419) );
  NAND2XL U2472 ( .A(n2456), .B(n2711), .Y(n2534) );
  NAND2XL U2473 ( .A(col[0]), .B(col[2]), .Y(n2193) );
  NAND2XL U2474 ( .A(col[2]), .B(n2672), .Y(n2208) );
  OR2XL U2475 ( .A(n2534), .B(n2070), .Y(n2071) );
  NAND2XL U2476 ( .A(n2711), .B(col[1]), .Y(n2181) );
  NAND2XL U2477 ( .A(n2170), .B(n2532), .Y(n2537) );
  NAND2XL U2478 ( .A(n2672), .B(n2455), .Y(n2222) );
  NAND2XL U2479 ( .A(n2174), .B(n2532), .Y(n2066) );
  AOI2BB1XL U2480 ( .A0N(n3007), .A1N(count_receive[1]), .B0(n2067), .Y(n2072)
         );
  NOR2X1 U2481 ( .A(n2068), .B(n2070), .Y(n2069) );
  INVXL U2482 ( .A(n2532), .Y(n2070) );
  NOR2X1 U2483 ( .A(count_out[2]), .B(n2975), .Y(n2529) );
  AOI2BB2XL U2484 ( .B0(n3082), .B1(n3081), .A0N(row_store[3]), .A1N(n3082), 
        .Y(n1392) );
  AOI2BB2XL U2485 ( .B0(n3082), .B1(n3080), .A0N(row_store[2]), .A1N(n3082), 
        .Y(n1393) );
  AOI2BB2XL U2486 ( .B0(n3082), .B1(n3079), .A0N(row_store[1]), .A1N(n3082), 
        .Y(n1394) );
  AOI2BB2XL U2487 ( .B0(n3082), .B1(n3078), .A0N(row_store[0]), .A1N(n3082), 
        .Y(n1395) );
  OAI21XL U2488 ( .A0(n2822), .A1(n2394), .B0(n2393), .Y(n1402) );
  NAND2XL U2489 ( .A(n2394), .B(y_array[6]), .Y(n2393) );
  AOI211XL U2490 ( .A0(row[1]), .A1(n2420), .B0(n2392), .C0(n2391), .Y(n2394)
         );
  OAI21XL U2491 ( .A0(n2822), .A1(n2409), .B0(n2408), .Y(n1406) );
  NAND2XL U2492 ( .A(n2409), .B(y_array[2]), .Y(n2408) );
  AOI211XL U2493 ( .A0(n2407), .A1(n2406), .B0(n2405), .C0(n2404), .Y(n2409)
         );
  OAI21XL U2494 ( .A0(n2822), .A1(n2387), .B0(n2386), .Y(n1407) );
  NAND2XL U2495 ( .A(n2387), .B(y_array[3]), .Y(n2386) );
  AOI211XL U2496 ( .A0(n2407), .A1(n2385), .B0(n2384), .C0(n2383), .Y(n2387)
         );
  OAI21XL U2497 ( .A0(n2822), .A1(n2375), .B0(n2374), .Y(n1454) );
  NAND2XL U2498 ( .A(n2375), .B(y_array[8]), .Y(n2374) );
  AOI211XL U2499 ( .A0(n2400), .A1(n2380), .B0(n2373), .C0(n2372), .Y(n2375)
         );
  NOR2X1 U2500 ( .A(n2371), .B(n2376), .Y(n2373) );
  OAI21XL U2501 ( .A0(n2822), .A1(n2382), .B0(n2381), .Y(n1456) );
  NAND2XL U2502 ( .A(n2382), .B(y_array[10]), .Y(n2381) );
  AOI211XL U2503 ( .A0(n2407), .A1(n2380), .B0(n2379), .C0(n2378), .Y(n2382)
         );
  OAI21XL U2504 ( .A0(n2822), .A1(n2365), .B0(n2364), .Y(n1455) );
  NAND2XL U2505 ( .A(n2365), .B(y_array[9]), .Y(n2364) );
  AOI211XL U2506 ( .A0(n2363), .A1(n2400), .B0(n2362), .C0(n2361), .Y(n2365)
         );
  NOR2X1 U2507 ( .A(n2371), .B(n2360), .Y(n2361) );
  OAI21XL U2508 ( .A0(n2822), .A1(n2354), .B0(n2353), .Y(n1457) );
  NAND2XL U2509 ( .A(n2354), .B(y_array[11]), .Y(n2353) );
  AOI211XL U2510 ( .A0(n2407), .A1(n2363), .B0(n2352), .C0(n2351), .Y(n2354)
         );
  OAI21XL U2511 ( .A0(n2822), .A1(n2369), .B0(n2368), .Y(n1405) );
  NAND2XL U2512 ( .A(n2369), .B(y_array[1]), .Y(n2368) );
  AOI211XL U2513 ( .A0(n2385), .A1(n2400), .B0(n2367), .C0(n2366), .Y(n2369)
         );
  OAI22XL U2514 ( .A0(n2502), .A1(n2515), .B0(n2517), .B1(n2568), .Y(n1474) );
  OAI2BB2XL U2515 ( .B0(n2577), .B1(n2568), .A0N(array_look_back[77]), .A1N(
        n2576), .Y(n1475) );
  OAI22XL U2516 ( .A0(n2438), .A1(n2568), .B0(n2437), .B1(n2436), .Y(n1476) );
  OAI2BB2XL U2517 ( .B0(n2575), .B1(n2568), .A0N(array_look_back[53]), .A1N(
        n2574), .Y(n1477) );
  OAI2BB2XL U2518 ( .B0(n2573), .B1(n2568), .A0N(array_look_back[41]), .A1N(
        n2572), .Y(n1478) );
  OAI2BB2XL U2519 ( .B0(n2571), .B1(n2568), .A0N(array_look_back[29]), .A1N(
        n2570), .Y(n1479) );
  OAI22XL U2520 ( .A0(n2504), .A1(n2515), .B0(n2517), .B1(n2560), .Y(n1522) );
  OAI2BB2XL U2521 ( .B0(n2577), .B1(n2560), .A0N(array_look_back[73]), .A1N(
        n2576), .Y(n1523) );
  OAI22XL U2522 ( .A0(n2438), .A1(n2560), .B0(n2432), .B1(n2436), .Y(n1524) );
  OAI2BB2XL U2523 ( .B0(n2575), .B1(n2560), .A0N(array_look_back[49]), .A1N(
        n2574), .Y(n1525) );
  OAI2BB2XL U2524 ( .B0(n2573), .B1(n2560), .A0N(array_look_back[37]), .A1N(
        n2572), .Y(n1526) );
  OAI2BB2XL U2525 ( .B0(n2571), .B1(n2560), .A0N(array_look_back[25]), .A1N(
        n2570), .Y(n1527) );
  OAI22XL U2526 ( .A0(n2517), .A1(n2562), .B0(n2514), .B1(n2515), .Y(n1510) );
  OAI2BB2XL U2527 ( .B0(n2577), .B1(n2562), .A0N(array_look_back[72]), .A1N(
        n2576), .Y(n1511) );
  OAI22XL U2528 ( .A0(n2438), .A1(n2562), .B0(n2429), .B1(n2436), .Y(n1512) );
  OAI2BB2XL U2529 ( .B0(n2575), .B1(n2562), .A0N(array_look_back[48]), .A1N(
        n2574), .Y(n1513) );
  OAI2BB2XL U2530 ( .B0(n2580), .B1(n2567), .A0N(n2578), .A1N(
        array_look_back[102]), .Y(n1485) );
  OAI22XL U2531 ( .A0(n2505), .A1(n2515), .B0(n2517), .B1(n2567), .Y(n1486) );
  OAI22XL U2532 ( .A0(n2577), .A1(n2567), .B0(n2909), .B1(n2499), .Y(n1487) );
  OAI22XL U2533 ( .A0(n2438), .A1(n2567), .B0(n2434), .B1(n2436), .Y(n1488) );
  OAI2BB2XL U2534 ( .B0(n2575), .B1(n2567), .A0N(array_look_back[54]), .A1N(
        n2574), .Y(n1489) );
  OAI2BB2XL U2535 ( .B0(n2566), .B1(n2567), .A0N(n2565), .A1N(
        array_look_back[18]), .Y(n1492) );
  OAI2BB2XL U2536 ( .B0(n2569), .B1(n2567), .A0N(n2792), .A1N(
        array_look_back[6]), .Y(n1493) );
  OAI22XL U2537 ( .A0(n2517), .A1(n2558), .B0(n2516), .B1(n2515), .Y(n1546) );
  OAI22XL U2538 ( .A0(n2577), .A1(n2558), .B0(n2955), .B1(n2499), .Y(n1547) );
  OAI22XL U2539 ( .A0(n2438), .A1(n2558), .B0(n2433), .B1(n2436), .Y(n1548) );
  OAI2BB2XL U2540 ( .B0(n2575), .B1(n2558), .A0N(array_look_back[51]), .A1N(
        n2574), .Y(n1549) );
  OAI2BB2XL U2541 ( .B0(n2580), .B1(n2556), .A0N(n2578), .A1N(
        array_look_back[107]), .Y(n1565) );
  OAI22XL U2542 ( .A0(n2506), .A1(n2515), .B0(n2517), .B1(n2556), .Y(n1569) );
  OAI2BB2XL U2543 ( .B0(n2577), .B1(n2556), .A0N(array_look_back[83]), .A1N(
        n2576), .Y(n1573) );
  OAI22XL U2544 ( .A0(n2438), .A1(n2556), .B0(n2428), .B1(n2436), .Y(n1577) );
  OAI2BB2XL U2545 ( .B0(n2575), .B1(n2556), .A0N(array_look_back[59]), .A1N(
        n2574), .Y(n1581) );
  OAI2BB2XL U2546 ( .B0(n2573), .B1(n2556), .A0N(array_look_back[47]), .A1N(
        n2572), .Y(n1585) );
  OAI2BB2XL U2547 ( .B0(n2571), .B1(n2556), .A0N(array_look_back[35]), .A1N(
        n2570), .Y(n1589) );
  OAI2BB2XL U2548 ( .B0(n2569), .B1(n2556), .A0N(n2792), .A1N(
        array_look_back[11]), .Y(n1597) );
  OAI22XL U2549 ( .A0(n2517), .A1(n2559), .B0(n2513), .B1(n2515), .Y(n1534) );
  OAI2BB2XL U2550 ( .B0(n2577), .B1(n2559), .A0N(array_look_back[74]), .A1N(
        n2576), .Y(n1535) );
  OAI22XL U2551 ( .A0(n2438), .A1(n2559), .B0(n2435), .B1(n2436), .Y(n1536) );
  OAI2BB2XL U2552 ( .B0(n2575), .B1(n2559), .A0N(array_look_back[50]), .A1N(
        n2574), .Y(n1537) );
  OAI2BB2XL U2553 ( .B0(n2573), .B1(n2559), .A0N(array_look_back[38]), .A1N(
        n2572), .Y(n1538) );
  OAI22XL U2554 ( .A0(n2501), .A1(n2515), .B0(n2517), .B1(n2557), .Y(n1570) );
  OAI22XL U2555 ( .A0(n2577), .A1(n2557), .B0(n2858), .B1(n2499), .Y(n1574) );
  OAI22XL U2556 ( .A0(n2438), .A1(n2557), .B0(n2430), .B1(n2436), .Y(n1578) );
  OAI2BB2XL U2557 ( .B0(n2575), .B1(n2557), .A0N(array_look_back[58]), .A1N(
        n2574), .Y(n1582) );
  OAI2BB2XL U2558 ( .B0(n2573), .B1(n2557), .A0N(array_look_back[46]), .A1N(
        n2572), .Y(n1586) );
  OAI22XL U2559 ( .A0(n2899), .A1(n2515), .B0(n2517), .B1(n2554), .Y(n1572) );
  OAI22XL U2560 ( .A0(n2891), .A1(n2499), .B0(n2577), .B1(n2554), .Y(n1576) );
  OAI22XL U2561 ( .A0(n2890), .A1(n2436), .B0(n2438), .B1(n2554), .Y(n1580) );
  OAI2BB2XL U2562 ( .B0(n2575), .B1(n2554), .A0N(array_look_back[56]), .A1N(
        n2574), .Y(n1584) );
  OAI2BB2XL U2563 ( .B0(n2571), .B1(n2554), .A0N(array_look_back[32]), .A1N(
        n2570), .Y(n1592) );
  OAI22XL U2564 ( .A0(n2503), .A1(n2515), .B0(n2517), .B1(n2555), .Y(n1571) );
  OAI2BB2XL U2565 ( .B0(n2577), .B1(n2555), .A0N(array_look_back[81]), .A1N(
        n2576), .Y(n1575) );
  OAI22XL U2566 ( .A0(n2427), .A1(n2436), .B0(n2438), .B1(n2555), .Y(n1579) );
  OAI2BB2XL U2567 ( .B0(n2575), .B1(n2555), .A0N(array_look_back[57]), .A1N(
        n2574), .Y(n1583) );
  OAI2BB2XL U2568 ( .B0(n2573), .B1(n2555), .A0N(array_look_back[45]), .A1N(
        n2572), .Y(n1587) );
  OAI2BB2XL U2569 ( .B0(n2571), .B1(n2555), .A0N(array_look_back[33]), .A1N(
        n2570), .Y(n1591) );
  OAI21XL U2570 ( .A0(n2822), .A1(n2359), .B0(n2358), .Y(n1403) );
  NAND2XL U2571 ( .A(n2359), .B(y_array[7]), .Y(n2358) );
  OAI22XL U2572 ( .A0(n2390), .A1(n2410), .B0(n3079), .B1(n2411), .Y(n2356) );
  OAI22XL U2573 ( .A0(n2846), .A1(n2515), .B0(n2517), .B1(n2564), .Y(n1498) );
  OAI22XL U2574 ( .A0(n2577), .A1(n2564), .B0(n2843), .B1(n2499), .Y(n1499) );
  OAI22XL U2575 ( .A0(n2438), .A1(n2564), .B0(n2845), .B1(n2436), .Y(n1500) );
  OAI2BB2XL U2576 ( .B0(n2575), .B1(n2564), .A0N(array_look_back[55]), .A1N(
        n2574), .Y(n1501) );
  OAI2BB2XL U2577 ( .B0(n2573), .B1(n2564), .A0N(array_look_back[43]), .A1N(
        n2572), .Y(n1502) );
  OAI21XL U2578 ( .A0(n2822), .A1(n2402), .B0(n2401), .Y(n1404) );
  NAND2XL U2579 ( .A(n2402), .B(y_array[0]), .Y(n2401) );
  AOI211XL U2580 ( .A0(n2406), .A1(n2400), .B0(n2399), .C0(n2398), .Y(n2402)
         );
  OAI22XL U2581 ( .A0(n2500), .A1(n2515), .B0(n2517), .B1(n2579), .Y(n1462) );
  OAI2BB2XL U2582 ( .B0(n2577), .B1(n2579), .A0N(array_look_back[76]), .A1N(
        n2576), .Y(n1463) );
  OAI22XL U2583 ( .A0(n2438), .A1(n2579), .B0(n2431), .B1(n2436), .Y(n1464) );
  OAI2BB2XL U2584 ( .B0(n2575), .B1(n2579), .A0N(array_look_back[52]), .A1N(
        n2574), .Y(n1465) );
  OAI2BB2XL U2585 ( .B0(n2573), .B1(n2579), .A0N(array_look_back[40]), .A1N(
        n2572), .Y(n1466) );
  OAI2BB2XL U2586 ( .B0(n2571), .B1(n2579), .A0N(array_look_back[28]), .A1N(
        n2570), .Y(n1467) );
  OAI21XL U2587 ( .A0(n2822), .A1(n2415), .B0(n2414), .Y(n1401) );
  NAND2XL U2588 ( .A(n2415), .B(y_array[5]), .Y(n2414) );
  OAI22XL U2589 ( .A0(row[1]), .A1(n2411), .B0(n2417), .B1(n2410), .Y(n2412)
         );
  MXI2XL U2590 ( .A(n2822), .B(n2803), .S0(n2802), .Y(n1411) );
  MXI2XL U2591 ( .A(n2822), .B(n2791), .S0(n2790), .Y(n1412) );
  INVXL U2592 ( .A(n2785), .Y(n2786) );
  MXI2XL U2593 ( .A(n2780), .B(n2822), .S0(n2779), .Y(n1413) );
  MXI2XL U2594 ( .A(n2822), .B(n2773), .S0(n2772), .Y(n1414) );
  MXI2XL U2595 ( .A(n2822), .B(n2753), .S0(n2752), .Y(n1416) );
  MXI2XL U2596 ( .A(n2822), .B(n2743), .S0(n2742), .Y(n1419) );
  MXI2XL U2597 ( .A(n2822), .B(n2738), .S0(n2737), .Y(n1420) );
  MXI2XL U2598 ( .A(n2822), .B(n2724), .S0(n2723), .Y(n1424) );
  MXI2XL U2599 ( .A(n2822), .B(n2720), .S0(n2719), .Y(n1426) );
  OAI22XL U2600 ( .A0(n2512), .A1(n3007), .B0(n2511), .B1(n2822), .Y(n1431) );
  NAND2XL U2601 ( .A(n2511), .B(sub_array[10]), .Y(n2512) );
  OAI22XL U2602 ( .A0(n2509), .A1(n3007), .B0(n2508), .B1(n2822), .Y(n1432) );
  NAND2XL U2603 ( .A(n2508), .B(sub_array[8]), .Y(n2509) );
  AOI222XL U2604 ( .A0(n2507), .A1(n2510), .B0(n2629), .B1(n2650), .C0(n2652), 
        .C1(n2628), .Y(n2508) );
  OAI22XL U2605 ( .A0(n2478), .A1(n3007), .B0(n2477), .B1(n2822), .Y(n1433) );
  NAND2XL U2606 ( .A(n2477), .B(sub_array[2]), .Y(n2478) );
  AOI222XL U2607 ( .A0(n2518), .A1(n2476), .B0(n2620), .B1(n2645), .C0(n2623), 
        .C1(n2644), .Y(n2477) );
  OAI22XL U2608 ( .A0(n2474), .A1(n3007), .B0(n2473), .B1(n2822), .Y(n1434) );
  NAND2XL U2609 ( .A(n2473), .B(sub_array[0]), .Y(n2474) );
  AOI222XL U2610 ( .A0(n2507), .A1(n2476), .B0(n2629), .B1(n2644), .C0(n2645), 
        .C1(n2628), .Y(n2473) );
  MXI2XL U2611 ( .A(n2658), .B(n2822), .S0(n2657), .Y(n1435) );
  OAI211XL U2612 ( .A0(n2656), .A1(n2655), .B0(n2654), .C0(n2792), .Y(n2657)
         );
  AOI22XL U2613 ( .A0(n2653), .A1(n2652), .B0(n2651), .B1(n2650), .Y(n2654) );
  MXI2XL U2614 ( .A(n2649), .B(n2822), .S0(n2648), .Y(n1436) );
  OAI211XL U2615 ( .A0(n2656), .A1(n2647), .B0(n2646), .C0(n2792), .Y(n2648)
         );
  AOI22XL U2616 ( .A0(n2653), .A1(n2645), .B0(n2651), .B1(n2644), .Y(n2646) );
  OAI21XL U2617 ( .A0(n2822), .A1(n2488), .B0(n2487), .Y(n1437) );
  NAND2XL U2618 ( .A(n2488), .B(sub_array[7]), .Y(n2487) );
  AOI211XL U2619 ( .A0(n2611), .A1(n2652), .B0(n3007), .C0(n2486), .Y(n2488)
         );
  OAI22XL U2620 ( .A0(n2490), .A1(n2655), .B0(n2592), .B1(n2485), .Y(n2486) );
  OAI21XL U2621 ( .A0(n2822), .A1(n2525), .B0(n2524), .Y(n1438) );
  NAND2XL U2622 ( .A(n2525), .B(sub_array[6]), .Y(n2524) );
  MXI2XL U2623 ( .A(n2822), .B(n2643), .S0(n2642), .Y(n1439) );
  AOI222XL U2624 ( .A0(n2641), .A1(n2640), .B0(n2651), .B1(n2639), .C0(n2638), 
        .C1(n2653), .Y(n2642) );
  OAI21XL U2625 ( .A0(n2822), .A1(n2521), .B0(n2520), .Y(n1440) );
  NAND2XL U2626 ( .A(n2521), .B(sub_array[4]), .Y(n2520) );
  AOI222XL U2627 ( .A0(n2641), .A1(n2630), .B0(n2629), .B1(n2639), .C0(n2638), 
        .C1(n2628), .Y(n2521) );
  OAI21XL U2628 ( .A0(n2822), .A1(n2523), .B0(n2522), .Y(n1441) );
  NAND2XL U2629 ( .A(n2523), .B(sub_array[3]), .Y(n2522) );
  AOI222XL U2630 ( .A0(n2641), .A1(n2613), .B0(n2612), .B1(n2639), .C0(n2638), 
        .C1(n2611), .Y(n2523) );
  OAI21XL U2631 ( .A0(n2822), .A1(n2498), .B0(n2497), .Y(n1442) );
  NAND2XL U2632 ( .A(n2498), .B(sub_array[22]), .Y(n2497) );
  AOI222XL U2633 ( .A0(n2635), .A1(n2624), .B0(n2623), .B1(n2634), .C0(n2633), 
        .C1(n2620), .Y(n2498) );
  MXI2XL U2634 ( .A(n2822), .B(n2637), .S0(n2636), .Y(n1443) );
  AOI222XL U2635 ( .A0(n2635), .A1(n2640), .B0(n2651), .B1(n2634), .C0(n2633), 
        .C1(n2653), .Y(n2636) );
  MXI2XL U2636 ( .A(n2822), .B(n2632), .S0(n2631), .Y(n1444) );
  AOI222XL U2637 ( .A0(n2635), .A1(n2630), .B0(n2629), .B1(n2634), .C0(n2633), 
        .C1(n2628), .Y(n2631) );
  OAI21XL U2638 ( .A0(n2822), .A1(n2496), .B0(n2495), .Y(n1445) );
  NAND2XL U2639 ( .A(n2496), .B(sub_array[19]), .Y(n2495) );
  AOI222XL U2640 ( .A0(n2635), .A1(n2613), .B0(n2612), .B1(n2634), .C0(n2633), 
        .C1(n2611), .Y(n2496) );
  MXI2XL U2641 ( .A(n2822), .B(n2627), .S0(n2626), .Y(n1446) );
  MXI2XL U2642 ( .A(n2822), .B(n2619), .S0(n2618), .Y(n1447) );
  AOI222XL U2643 ( .A0(n2625), .A1(n2640), .B0(n2651), .B1(n2622), .C0(n2621), 
        .C1(n2653), .Y(n2618) );
  MXI2XL U2644 ( .A(n2822), .B(n2617), .S0(n2616), .Y(n1448) );
  AOI222XL U2645 ( .A0(n2625), .A1(n2630), .B0(n2629), .B1(n2622), .C0(n2621), 
        .C1(n2628), .Y(n2616) );
  MXI2XL U2646 ( .A(n2822), .B(n2615), .S0(n2614), .Y(n1449) );
  AOI222XL U2647 ( .A0(n2625), .A1(n2613), .B0(n2612), .B1(n2622), .C0(n2621), 
        .C1(n2611), .Y(n2614) );
  MXI2XL U2648 ( .A(n2822), .B(n2601), .S0(n2600), .Y(n1450) );
  AOI222XL U2649 ( .A0(n2624), .A1(n2599), .B0(n2598), .B1(n2623), .C0(n2620), 
        .C1(n2597), .Y(n2600) );
  MXI2XL U2650 ( .A(n2822), .B(n2596), .S0(n2595), .Y(n1451) );
  AOI222XL U2651 ( .A0(n2640), .A1(n2599), .B0(n2598), .B1(n2651), .C0(n2653), 
        .C1(n2597), .Y(n2595) );
  MXI2XL U2652 ( .A(n2822), .B(n2590), .S0(n2589), .Y(n1452) );
  AOI222XL U2653 ( .A0(n2630), .A1(n2599), .B0(n2598), .B1(n2629), .C0(n2628), 
        .C1(n2597), .Y(n2589) );
  MXI2XL U2654 ( .A(n2822), .B(n2588), .S0(n2587), .Y(n1453) );
  AOI222XL U2655 ( .A0(n2599), .A1(n2613), .B0(n2611), .B1(n2597), .C0(n2612), 
        .C1(n2598), .Y(n2587) );
  AOI21XL U2656 ( .A0(n2314), .A1(n2425), .B0(n2223), .Y(n2225) );
  AOI211XL U2657 ( .A0(n2425), .A1(n2313), .B0(n2213), .C0(n2539), .Y(n2215)
         );
  AOI211XL U2658 ( .A0(n2425), .A1(n2311), .B0(n2175), .C0(n2540), .Y(n2177)
         );
  AOI211XL U2659 ( .A0(n2425), .A1(n2303), .B0(n2182), .C0(n2541), .Y(n2184)
         );
  AOI211XL U2660 ( .A0(n2425), .A1(n2306), .B0(n2209), .C0(n2542), .Y(n2211)
         );
  AOI211XL U2661 ( .A0(n2425), .A1(n2305), .B0(n2194), .C0(n2543), .Y(n2196)
         );
  AOI211XL U2662 ( .A0(n2425), .A1(n2310), .B0(n2199), .C0(n2544), .Y(n2201)
         );
  AOI211XL U2663 ( .A0(n2425), .A1(n2309), .B0(n2185), .C0(n2545), .Y(n2187)
         );
  AOI211XL U2664 ( .A0(n2425), .A1(n2312), .B0(n2189), .C0(n2546), .Y(n2191)
         );
  AOI211XL U2665 ( .A0(n2425), .A1(n2308), .B0(n2217), .C0(n2547), .Y(n2219)
         );
  AOI211XL U2666 ( .A0(n2425), .A1(n2307), .B0(n2204), .C0(n2548), .Y(n2206)
         );
  AOI2BB2XL U2667 ( .B0(n2551), .B1(n2552), .A0N(n2552), .A1N(row_store[46]), 
        .Y(n1617) );
  AOI2BB2XL U2668 ( .B0(n2551), .B1(n2548), .A0N(n2548), .A1N(row_store[42]), 
        .Y(n1621) );
  AOI2BB2XL U2669 ( .B0(n2551), .B1(n2547), .A0N(n2547), .A1N(row_store[38]), 
        .Y(n1625) );
  AOI2BB2XL U2670 ( .B0(n2551), .B1(n2546), .A0N(n2546), .A1N(row_store[34]), 
        .Y(n1629) );
  AOI2BB2XL U2671 ( .B0(n2551), .B1(n2545), .A0N(n2545), .A1N(row_store[30]), 
        .Y(n1633) );
  AOI2BB2XL U2672 ( .B0(n2551), .B1(n2544), .A0N(n2544), .A1N(row_store[26]), 
        .Y(n1637) );
  AOI2BB2XL U2673 ( .B0(n2551), .B1(n2543), .A0N(n2543), .A1N(row_store[22]), 
        .Y(n1641) );
  AOI2BB2XL U2674 ( .B0(n2551), .B1(n2542), .A0N(n2542), .A1N(row_store[18]), 
        .Y(n1645) );
  AOI2BB2XL U2675 ( .B0(n2551), .B1(n2541), .A0N(n2541), .A1N(row_store[14]), 
        .Y(n1649) );
  AOI2BB2XL U2676 ( .B0(n2551), .B1(n2540), .A0N(n2540), .A1N(row_store[10]), 
        .Y(n1653) );
  AOI2BB2XL U2677 ( .B0(n2551), .B1(n2539), .A0N(n2539), .A1N(row_store[6]), 
        .Y(n1657) );
  AOI2BB2XL U2678 ( .B0(n2549), .B1(n2552), .A0N(n2552), .A1N(row_store[44]), 
        .Y(n1619) );
  AOI2BB2XL U2679 ( .B0(n2549), .B1(n2548), .A0N(n2548), .A1N(row_store[40]), 
        .Y(n1623) );
  AOI2BB2XL U2680 ( .B0(n2549), .B1(n2547), .A0N(n2547), .A1N(row_store[36]), 
        .Y(n1627) );
  AOI2BB2XL U2681 ( .B0(n2549), .B1(n2546), .A0N(n2546), .A1N(row_store[32]), 
        .Y(n1631) );
  AOI2BB2XL U2682 ( .B0(n2549), .B1(n2545), .A0N(n2545), .A1N(row_store[28]), 
        .Y(n1635) );
  AOI2BB2XL U2683 ( .B0(n2549), .B1(n2544), .A0N(n2544), .A1N(row_store[24]), 
        .Y(n1639) );
  AOI2BB2XL U2684 ( .B0(n2549), .B1(n2543), .A0N(n2543), .A1N(row_store[20]), 
        .Y(n1643) );
  AOI2BB2XL U2685 ( .B0(n2549), .B1(n2542), .A0N(n2542), .A1N(row_store[16]), 
        .Y(n1647) );
  AOI2BB2XL U2686 ( .B0(n2549), .B1(n2541), .A0N(n2541), .A1N(row_store[12]), 
        .Y(n1651) );
  AOI2BB2XL U2687 ( .B0(n2549), .B1(n2540), .A0N(n2540), .A1N(row_store[8]), 
        .Y(n1655) );
  AOI2BB2XL U2688 ( .B0(n2549), .B1(n2539), .A0N(n2539), .A1N(row_store[4]), 
        .Y(n1659) );
  AOI2BB2XL U2689 ( .B0(n2550), .B1(n2552), .A0N(n2552), .A1N(row_store[47]), 
        .Y(n1618) );
  AOI2BB2XL U2690 ( .B0(n2550), .B1(n2548), .A0N(n2548), .A1N(row_store[43]), 
        .Y(n1622) );
  AOI2BB2XL U2691 ( .B0(n2550), .B1(n2547), .A0N(n2547), .A1N(row_store[39]), 
        .Y(n1626) );
  AOI2BB2XL U2692 ( .B0(n2550), .B1(n2546), .A0N(n2546), .A1N(row_store[35]), 
        .Y(n1630) );
  AOI2BB2XL U2693 ( .B0(n2550), .B1(n2545), .A0N(n2545), .A1N(row_store[31]), 
        .Y(n1634) );
  AOI2BB2XL U2694 ( .B0(n2550), .B1(n2544), .A0N(n2544), .A1N(row_store[27]), 
        .Y(n1638) );
  AOI2BB2XL U2695 ( .B0(n2550), .B1(n2543), .A0N(n2543), .A1N(row_store[23]), 
        .Y(n1642) );
  AOI2BB2XL U2696 ( .B0(n2550), .B1(n2542), .A0N(n2542), .A1N(row_store[19]), 
        .Y(n1646) );
  AOI2BB2XL U2697 ( .B0(n2550), .B1(n2541), .A0N(n2541), .A1N(row_store[15]), 
        .Y(n1650) );
  AOI2BB2XL U2698 ( .B0(n2550), .B1(n2540), .A0N(n2540), .A1N(row_store[11]), 
        .Y(n1654) );
  AOI2BB2XL U2699 ( .B0(n2550), .B1(n2539), .A0N(n2539), .A1N(row_store[7]), 
        .Y(n1658) );
  AOI2BB2XL U2700 ( .B0(n2553), .B1(n2539), .A0N(n2539), .A1N(row_store[5]), 
        .Y(n1656) );
  AOI2BB2XL U2701 ( .B0(n2553), .B1(n2541), .A0N(n2541), .A1N(row_store[13]), 
        .Y(n1648) );
  AOI2BB2XL U2702 ( .B0(n2553), .B1(n2547), .A0N(n2547), .A1N(row_store[37]), 
        .Y(n1624) );
  AOI2BB2XL U2703 ( .B0(n2553), .B1(n2552), .A0N(n2552), .A1N(row_store[45]), 
        .Y(n1616) );
  AOI2BB2XL U2704 ( .B0(n2553), .B1(n2540), .A0N(n2540), .A1N(row_store[9]), 
        .Y(n1652) );
  AOI2BB2XL U2705 ( .B0(n2553), .B1(n2544), .A0N(n2544), .A1N(row_store[25]), 
        .Y(n1636) );
  AOI2BB2XL U2706 ( .B0(n2553), .B1(n2542), .A0N(n2542), .A1N(row_store[17]), 
        .Y(n1644) );
  AOI2BB2XL U2707 ( .B0(n2553), .B1(n2543), .A0N(n2543), .A1N(row_store[21]), 
        .Y(n1640) );
  AOI2BB2XL U2708 ( .B0(n2553), .B1(n2545), .A0N(n2545), .A1N(row_store[29]), 
        .Y(n1632) );
  AOI2BB2XL U2709 ( .B0(n2553), .B1(n2546), .A0N(n2546), .A1N(row_store[33]), 
        .Y(n1628) );
  AOI2BB2XL U2710 ( .B0(n2553), .B1(n2548), .A0N(n2548), .A1N(row_store[41]), 
        .Y(n1620) );
  AOI221XL U2711 ( .A0(n2529), .A1(current_state[2]), .B0(n1691), .B1(
        current_state[2]), .C0(n1690), .Y(n1685) );
  NOR2X1 U2712 ( .A(n2080), .B(n2079), .Y(n2082) );
  OAI2BB1XL U2713 ( .A0N(n2039), .A1N(n2987), .B0(n2038), .Y(n2051) );
  OAI21XL U2714 ( .A0(n2822), .A1(n2422), .B0(n2421), .Y(n1400) );
  NAND2XL U2715 ( .A(n2422), .B(y_array[4]), .Y(n2421) );
  AOI211XL U2716 ( .A0(n2420), .A1(n3079), .B0(n2419), .C0(n2418), .Y(n2422)
         );
  OAI2BB2XL U2717 ( .B0(col[1]), .B1(n2535), .A0N(n2792), .A1N(array_in[8]), 
        .Y(n1667) );
  NOR2X2 U2718 ( .A(n2697), .B(n2699), .Y(n2822) );
  AND2X2 U2719 ( .A(n2107), .B(n2032), .Y(n2307) );
  INVX2 U2720 ( .A(n2446), .Y(n2207) );
  INVXL U2721 ( .A(n1960), .Y(n1783) );
  INVXL U2722 ( .A(n2079), .Y(n2030) );
  INVXL U2723 ( .A(n2797), .Y(n2718) );
  XOR2XL U2724 ( .A(n2669), .B(n2450), .Y(n2602) );
  NOR2X2 U2725 ( .A(n2471), .B(x[0]), .Y(n1987) );
  INVXL U2726 ( .A(row[1]), .Y(n3079) );
  INVXL U2727 ( .A(n2366), .Y(n2560) );
  AOI222XL U2728 ( .A0(n2518), .A1(n2510), .B0(n2620), .B1(n2652), .C0(n2623), 
        .C1(n2650), .Y(n2511) );
  AOI222XL U2729 ( .A0(n2641), .A1(n2624), .B0(n2623), .B1(n2639), .C0(n2638), 
        .C1(n2620), .Y(n2525) );
  AOI222XL U2730 ( .A0(n2625), .A1(n2624), .B0(n2623), .B1(n2622), .C0(n2621), 
        .C1(n2620), .Y(n2626) );
  NAND2XL U2731 ( .A(count_out[0]), .B(count_out[1]), .Y(n2526) );
  INVXL U2732 ( .A(count_out[3]), .Y(n2833) );
  INVXL U2733 ( .A(n3056), .Y(n2975) );
  INVXL U2734 ( .A(current_state[0]), .Y(n2024) );
  INVXL U2735 ( .A(n2046), .Y(n1691) );
  INVXL U2736 ( .A(current_state[2]), .Y(n1998) );
  INVXL U2737 ( .A(count_receive[3]), .Y(n2074) );
  OAI22XL U2738 ( .A0(count[3]), .A1(n2074), .B0(n3083), .B1(count_receive[0]), 
        .Y(n1686) );
  AOI221XL U2739 ( .A0(n2074), .A1(count[3]), .B0(n3083), .B1(count_receive[0]), .C0(n1686), .Y(n1689) );
  INVXL U2740 ( .A(count_receive[1]), .Y(n2003) );
  OAI22XL U2741 ( .A0(count[1]), .A1(n2003), .B0(n3084), .B1(count_receive[2]), 
        .Y(n1687) );
  AOI221XL U2742 ( .A0(n2003), .A1(count[1]), .B0(n3084), .B1(count_receive[2]), .C0(n1687), .Y(n1688) );
  NAND3BXL U2743 ( .AN(n2169), .B(n1689), .C(n1688), .Y(n1999) );
  INVXL U2744 ( .A(n1999), .Y(n1690) );
  NAND2XL U2745 ( .A(current_state[2]), .B(n2046), .Y(n3086) );
  INVXL U2746 ( .A(count_out[1]), .Y(n2827) );
  INVXL U2747 ( .A(n2526), .Y(n2832) );
  AOI211XL U2748 ( .A0(n3085), .A1(n2827), .B0(n2832), .C0(n3086), .Y(N6083)
         );
  NAND2XL U2749 ( .A(count_out[2]), .B(n2832), .Y(n1692) );
  NAND2XL U2750 ( .A(count_out[3]), .B(n1692), .Y(n1693) );
  INVXL U2751 ( .A(n3059), .Y(n2898) );
  AOI21XL U2752 ( .A0(n1693), .A1(n2898), .B0(n3086), .Y(N6085) );
  INVX1 U2753 ( .A(n1987), .Y(n1864) );
  OAI211XL U2754 ( .A0(array_in[11]), .A1(n2202), .B0(n2116), .C0(x[1]), .Y(
        n1997) );
  NAND2XL U2755 ( .A(array_in[10]), .B(array_in[11]), .Y(n2035) );
  NAND2X1 U2756 ( .A(n2018), .B(n1931), .Y(n2569) );
  AOI32XL U2757 ( .A0(n2119), .A1(array_in[2]), .A2(array_in[1]), .B0(n2149), 
        .B1(array_in[2]), .Y(n1694) );
  INVXL U2758 ( .A(array_in[3]), .Y(n2103) );
  AOI32XL U2759 ( .A0(n2571), .A1(n2573), .A2(n1694), .B0(n2103), .B1(n2573), 
        .Y(n1695) );
  AOI32XL U2760 ( .A0(array_in[4]), .A1(array_in[5]), .A2(n1695), .B0(n2424), 
        .B1(array_in[5]), .Y(n1696) );
  NAND2X2 U2761 ( .A(n1987), .B(n1958), .Y(n2577) );
  NAND2X1 U2762 ( .A(n1908), .B(n1958), .Y(n2438) );
  INVXL U2763 ( .A(array_in[6]), .Y(n2987) );
  AOI32XL U2764 ( .A0(n1696), .A1(n2577), .A2(n2438), .B0(n2987), .B1(n2577), 
        .Y(n1697) );
  INVXL U2765 ( .A(n2005), .Y(n1961) );
  INVXL U2766 ( .A(n2048), .Y(n1698) );
  AOI222XL U2767 ( .A0(n1699), .A1(n1698), .B0(n1970), .B1(array_in[9]), .C0(
        n1918), .C1(n2116), .Y(n1996) );
  AOI22XL U2768 ( .A0(n1972), .A1(array_look_back[115]), .B0(n1966), .B1(
        array_look_back[55]), .Y(n1719) );
  AOI22XL U2769 ( .A0(n1973), .A1(array_look_back[67]), .B0(n1961), .B1(
        array_look_back[91]), .Y(n1725) );
  AOI22XL U2770 ( .A0(n1972), .A1(array_look_back[114]), .B0(n1966), .B1(
        array_look_back[54]), .Y(n1740) );
  AOI22XL U2771 ( .A0(n1973), .A1(array_look_back[66]), .B0(n1961), .B1(
        array_look_back[90]), .Y(n1746) );
  AOI22XL U2772 ( .A0(n1972), .A1(array_look_back[112]), .B0(n1961), .B1(
        array_look_back[88]), .Y(n1777) );
  AOI222XL U2773 ( .A0(n2018), .A1(add_array[11]), .B0(n2116), .B1(
        add_array[19]), .C0(n1958), .C1(add_array[15]), .Y(n1848) );
  INVXL U2774 ( .A(sub_array[13]), .Y(n2596) );
  OAI21XL U2775 ( .A0(sub_array[9]), .A1(add_array[20]), .B0(n2116), .Y(n1793)
         );
  OAI21XL U2776 ( .A0(n2007), .A1(n2596), .B0(n1793), .Y(n1798) );
  AOI22XL U2777 ( .A0(add_array[22]), .A1(n2116), .B0(add_array[18]), .B1(
        n1958), .Y(n1796) );
  NAND2XL U2778 ( .A(n1867), .B(n1796), .Y(n1797) );
  AOI22XL U2779 ( .A0(n1967), .A1(array_look_back[131]), .B0(sub_array[4]), 
        .B1(n2424), .Y(n1809) );
  INVXL U2780 ( .A(add_array[12]), .Y(n2724) );
  INVXL U2781 ( .A(n2438), .Y(n2426) );
  AOI22XL U2782 ( .A0(n1966), .A1(array_look_back[59]), .B0(add_array[16]), 
        .B1(n2426), .Y(n1800) );
  OAI21XL U2783 ( .A0(add_array[13]), .A1(array_look_back[35]), .B0(n2167), 
        .Y(n1799) );
  INVXL U2784 ( .A(array_look_back[23]), .Y(n2869) );
  INVXL U2785 ( .A(sub_array[1]), .Y(n2649) );
  AOI21XL U2786 ( .A0(n2869), .A1(n2649), .B0(n2566), .Y(n1801) );
  AOI211XL U2787 ( .A0(array_look_back[119]), .A1(n1972), .B0(n1802), .C0(
        n1801), .Y(n1806) );
  AOI22XL U2788 ( .A0(n1973), .A1(array_look_back[71]), .B0(n1968), .B1(
        array_look_back[83]), .Y(n1805) );
  AOI22XL U2789 ( .A0(n1969), .A1(array_look_back[143]), .B0(sub_array[12]), 
        .B1(n1979), .Y(n1804) );
  OAI21XL U2790 ( .A0(add_array[14]), .A1(array_look_back[47]), .B0(n2179), 
        .Y(n1803) );
  INVXL U2791 ( .A(add_array[21]), .Y(n2791) );
  INVXL U2792 ( .A(add_array[17]), .Y(n2773) );
  AOI22XL U2793 ( .A0(n1967), .A1(array_look_back[128]), .B0(n1973), .B1(
        array_look_back[68]), .Y(n1823) );
  AOI22XL U2794 ( .A0(n1972), .A1(array_look_back[116]), .B0(n1971), .B1(
        array_look_back[104]), .Y(n1820) );
  INVXL U2795 ( .A(array_look_back[56]), .Y(n2902) );
  AOI22XL U2796 ( .A0(n1967), .A1(array_look_back[129]), .B0(n1969), .B1(
        array_look_back[141]), .Y(n1842) );
  AOI22XL U2797 ( .A0(n1966), .A1(array_look_back[57]), .B0(n1968), .B1(
        array_look_back[81]), .Y(n1841) );
  AOI22XL U2798 ( .A0(n1961), .A1(array_look_back[93]), .B0(n1971), .B1(
        array_look_back[105]), .Y(n1840) );
  AOI22XL U2799 ( .A0(n1973), .A1(array_look_back[69]), .B0(n1972), .B1(
        array_look_back[117]), .Y(n1839) );
  INVXL U2800 ( .A(array_look_back[9]), .Y(n2151) );
  AOI221XL U2801 ( .A0(add_array[12]), .A1(n2179), .B0(array_look_back[45]), 
        .B1(n2179), .C0(y_array[9]), .Y(n1843) );
  INVXL U2802 ( .A(add_array[16]), .Y(n2803) );
  NAND2XL U2803 ( .A(n2116), .B(add_array[20]), .Y(n1865) );
  INVXL U2804 ( .A(n1856), .Y(n1857) );
  AOI2BB1XL U2805 ( .A0N(sub_array[1]), .A1N(array_look_back[10]), .B0(n2569), 
        .Y(n1868) );
  AOI211XL U2806 ( .A0(array_look_back[130]), .A1(n1967), .B0(y_array[10]), 
        .C0(n1868), .Y(n1876) );
  AOI22XL U2807 ( .A0(n1972), .A1(array_look_back[118]), .B0(add_array[16]), 
        .B1(n2006), .Y(n1875) );
  AOI22XL U2808 ( .A0(n1966), .A1(array_look_back[58]), .B0(sub_array[9]), 
        .B1(n1970), .Y(n1874) );
  AOI22XL U2809 ( .A0(n1968), .A1(array_look_back[82]), .B0(sub_array[13]), 
        .B1(n1979), .Y(n1872) );
  AOI22XL U2810 ( .A0(n2167), .A1(add_array[12]), .B0(n1961), .B1(
        array_look_back[94]), .Y(n1871) );
  AOI22XL U2811 ( .A0(n1973), .A1(array_look_back[70]), .B0(sub_array[5]), 
        .B1(n2424), .Y(n1870) );
  AOI22XL U2812 ( .A0(n1969), .A1(array_look_back[142]), .B0(n1971), .B1(
        array_look_back[106]), .Y(n1869) );
  AOI222XL U2813 ( .A0(n2018), .A1(sub_array[11]), .B0(n2116), .B1(
        sub_array[19]), .C0(n1958), .C1(sub_array[15]), .Y(n1907) );
  INVXL U2814 ( .A(sub_array[20]), .Y(n2632) );
  AOI22XL U2815 ( .A0(n1887), .A1(add_array[14]), .B0(n2116), .B1(
        add_array[10]), .Y(n1888) );
  AOI221XL U2816 ( .A0(array_look_back[13]), .A1(n2149), .B0(add_array[2]), 
        .B1(n2149), .C0(y_array[1]), .Y(n1891) );
  INVXL U2817 ( .A(add_array[13]), .Y(n2753) );
  AOI22XL U2818 ( .A0(n1972), .A1(array_look_back[109]), .B0(n1969), .B1(
        array_look_back[133]), .Y(n1898) );
  AOI22XL U2819 ( .A0(n1967), .A1(array_look_back[121]), .B0(n1971), .B1(
        array_look_back[97]), .Y(n1896) );
  AOI222XL U2820 ( .A0(n1908), .A1(sub_array[20]), .B0(n1951), .B1(
        sub_array[22]), .C0(n1987), .C1(sub_array[21]), .Y(n1912) );
  NAND2X2 U2821 ( .A(n2464), .B(n1969), .Y(n2171) );
  INVXL U2822 ( .A(n2171), .Y(n2157) );
  INVXL U2823 ( .A(n2563), .Y(n2087) );
  INVXL U2824 ( .A(sub_array[16]), .Y(n2617) );
  INVXL U2825 ( .A(add_array[5]), .Y(n2738) );
  INVXL U2826 ( .A(add_array[8]), .Y(n2720) );
  INVXL U2827 ( .A(sub_array[17]), .Y(n2619) );
  INVXL U2828 ( .A(add_array[6]), .Y(n2710) );
  OAI2BB1XL U2829 ( .A0N(n2619), .A1N(n2710), .B0(n2006), .Y(n1916) );
  AOI22XL U2830 ( .A0(n1967), .A1(array_look_back[123]), .B0(n1969), .B1(
        array_look_back[135]), .Y(n1943) );
  AOI211XL U2831 ( .A0(n1997), .A1(n2035), .B0(n1996), .C0(n2025), .Y(n2527)
         );
  OR2XL U2832 ( .A(n2023), .B(current_state[0]), .Y(n2105) );
  OAI211XL U2833 ( .A0(n2527), .A1(n2023), .B0(n2105), .C0(n1999), .Y(n1684)
         );
  NAND2XL U2834 ( .A(in_valid_num), .B(in_num[0]), .Y(n2000) );
  NOR3X1 U2835 ( .A(current_state[2]), .B(current_state[1]), .C(
        current_state[0]), .Y(n3007) );
  INVX2 U2836 ( .A(n3007), .Y(n2792) );
  OAI211XL U2837 ( .A0(in_valid_num), .A1(n3083), .B0(n2000), .C0(n2792), .Y(
        n1663) );
  NAND2XL U2838 ( .A(in_valid_num), .B(in_num[2]), .Y(n2001) );
  OAI211XL U2839 ( .A0(in_valid_num), .A1(n3084), .B0(n2001), .C0(n2792), .Y(
        n1661) );
  INVXL U2840 ( .A(in_valid_num), .Y(n2538) );
  AOI22XL U2841 ( .A0(in_valid_num), .A1(in_num[1]), .B0(count[1]), .B1(n2538), 
        .Y(n2002) );
  NAND2XL U2842 ( .A(n2002), .B(n2792), .Y(n1660) );
  INVXL U2843 ( .A(count_receive[0]), .Y(n2068) );
  INVXL U2844 ( .A(n2067), .Y(n2530) );
  OAI32XL U2845 ( .A0(count_receive[1]), .A1(n2068), .A2(n2070), .B0(n2530), 
        .B1(n2003), .Y(n1678) );
  INVXL U2846 ( .A(array_in[9]), .Y(n2031) );
  NAND2XL U2847 ( .A(col[3]), .B(n2456), .Y(n2004) );
  OAI22XL U2848 ( .A0(n3007), .A1(n2031), .B0(n2537), .B1(n2004), .Y(n1666) );
  OAI22XL U2849 ( .A0(n3007), .A1(n2103), .B0(n2537), .B1(n2181), .Y(n1672) );
  INVXL U2850 ( .A(array_in[10]), .Y(n2107) );
  INVXL U2851 ( .A(array_in[2]), .Y(n2985) );
  INVXL U2852 ( .A(array_in[0]), .Y(n2533) );
  NOR2X2 U2853 ( .A(n2102), .B(n2012), .Y(n2304) );
  INVXL U2854 ( .A(array_in[7]), .Y(n2065) );
  INVXL U2855 ( .A(n2098), .Y(n2019) );
  INVX1 U2856 ( .A(n2662), .Y(n2192) );
  INVXL U2857 ( .A(array_in[5]), .Y(n2104) );
  INVXL U2858 ( .A(n2085), .Y(n2041) );
  NAND2XL U2859 ( .A(n2084), .B(n2041), .Y(n2028) );
  NAND2XL U2860 ( .A(n2029), .B(n2985), .Y(n2094) );
  OAI21XL U2861 ( .A0(array_in[3]), .A1(n2086), .B0(n2094), .Y(n2040) );
  NAND2XL U2862 ( .A(n2057), .B(n2063), .Y(n2079) );
  OAI21XL U2863 ( .A0(N4586), .A1(array_in[8]), .B0(n2030), .Y(n2088) );
  AOI31XL U2864 ( .A0(n2096), .A1(n2563), .A2(n2031), .B0(n2088), .Y(n2044) );
  NAND2XL U2865 ( .A(n2096), .B(n2107), .Y(n2089) );
  OAI211XL U2866 ( .A0(array_in[11]), .A1(n2032), .B0(n2044), .C0(n2089), .Y(
        n2033) );
  OAI31XL U2867 ( .A0(array_in[7]), .A1(n2078), .A2(n2079), .B0(n2033), .Y(
        n2037) );
  NAND2XL U2868 ( .A(array_in[1]), .B(array_in[0]), .Y(n2034) );
  NAND2XL U2869 ( .A(n2038), .B(n2052), .Y(n2059) );
  INVXL U2870 ( .A(array_in[4]), .Y(n2990) );
  NAND2XL U2871 ( .A(array_in[6]), .B(n2039), .Y(n2058) );
  OAI21XL U2872 ( .A0(n2048), .A1(n2035), .B0(array_in[7]), .Y(n2036) );
  AOI31XL U2873 ( .A0(n2042), .A1(n2084), .A2(n2041), .B0(n2040), .Y(n2043) );
  AOI2BB1XL U2874 ( .A0N(n2045), .A1N(n2044), .B0(n2692), .Y(n2050) );
  NAND2XL U2875 ( .A(array_in[7]), .B(n2047), .Y(n2109) );
  OAI22XL U2876 ( .A0(n2110), .A1(n2471), .B0(n2048), .B1(n2109), .Y(n2049) );
  AOI211XL U2877 ( .A0(n2052), .A1(n2051), .B0(n2050), .C0(n2049), .Y(n2053)
         );
  OAI211XL U2878 ( .A0(n2192), .A1(n2760), .B0(n2114), .C0(n2053), .Y(n1614)
         );
  OAI21XL U2879 ( .A0(n2056), .A1(n2055), .B0(n2054), .Y(n2446) );
  INVXL U2880 ( .A(n2057), .Y(n2062) );
  INVXL U2881 ( .A(n2058), .Y(n2060) );
  OAI22XL U2882 ( .A0(n2060), .A1(n2059), .B0(n2110), .B1(n2464), .Y(n2061) );
  AOI31XL U2883 ( .A0(n2699), .A1(n2063), .A2(n2062), .B0(n2061), .Y(n2064) );
  OAI211XL U2884 ( .A0(n2207), .A1(n2760), .B0(n2114), .C0(n2064), .Y(n1615)
         );
  NAND2XL U2885 ( .A(n2188), .B(n2532), .Y(n2535) );
  OAI22XL U2886 ( .A0(n3007), .A1(n2107), .B0(n2535), .B1(n2456), .Y(n1665) );
  OAI22XL U2887 ( .A0(n3007), .A1(n2987), .B0(n2066), .B1(n2208), .Y(n1669) );
  OAI22XL U2888 ( .A0(n3007), .A1(n2065), .B0(n2066), .B1(n2193), .Y(n1668) );
  OAI22XL U2889 ( .A0(n3007), .A1(n2985), .B0(n2066), .B1(n2222), .Y(n1673) );
  NAND2XL U2890 ( .A(count_receive[1]), .B(n2069), .Y(n2076) );
  INVXL U2891 ( .A(count_receive[2]), .Y(n2077) );
  AOI22XL U2892 ( .A0(count_receive[2]), .A1(n2072), .B0(n2076), .B1(n2077), 
        .Y(n1677) );
  OAI22XL U2893 ( .A0(n3007), .A1(n2990), .B0(n2071), .B1(n2208), .Y(n1671) );
  OAI22XL U2894 ( .A0(n3007), .A1(n2104), .B0(n2071), .B1(n2193), .Y(n1670) );
  OAI2BB1XL U2895 ( .A0N(n2077), .A1N(n2532), .B0(n2072), .Y(n2073) );
  INVXL U2896 ( .A(n2073), .Y(n2075) );
  OAI32XL U2897 ( .A0(count_receive[3]), .A1(n2077), .A2(n2076), .B0(n2075), 
        .B1(n2074), .Y(n1676) );
  INVXL U2898 ( .A(n2441), .Y(n2667) );
  AOI22XL U2899 ( .A0(n2699), .A1(n2082), .B0(n2425), .B1(n2667), .Y(n2083) );
  OAI211XL U2900 ( .A0(n2110), .A1(n2685), .B0(n2083), .C0(n2109), .Y(n1680)
         );
  OAI22XL U2901 ( .A0(array_in[3]), .A1(n2086), .B0(n2085), .B1(n2084), .Y(
        n2093) );
  AOI2BB1XL U2902 ( .A0N(n2090), .A1N(n2089), .B0(n2088), .Y(n2091) );
  AOI211XL U2903 ( .A0(n2094), .A1(n2093), .B0(n2092), .C0(n2091), .Y(n2115)
         );
  OAI211XL U2904 ( .A0(n2095), .A1(n2102), .B0(n2101), .C0(n2100), .Y(n2440)
         );
  AOI32XL U2905 ( .A0(array_in[4]), .A1(array_in[2]), .A2(n2104), .B0(n2103), 
        .B1(array_in[2]), .Y(n2106) );
  AOI211XL U2906 ( .A0(array_in[1]), .A1(n2106), .B0(n2533), .C0(n2105), .Y(
        n2112) );
  OAI22XL U2907 ( .A0(n2110), .A1(n2680), .B0(n2109), .B1(n2108), .Y(n2111) );
  AOI211XL U2908 ( .A0(n2425), .A1(n2440), .B0(n2112), .C0(n2111), .Y(n2113)
         );
  OAI211XL U2909 ( .A0(n2115), .A1(n2692), .B0(n2114), .C0(n2113), .Y(n1613)
         );
  INVXL U2910 ( .A(array_look_back[119]), .Y(n2870) );
  AOI221XL U2911 ( .A0(n2123), .A1(n2122), .B0(n2121), .B1(n2122), .C0(n2146), 
        .Y(n2125) );
  INVXL U2912 ( .A(n2126), .Y(n2142) );
  INVXL U2913 ( .A(n2127), .Y(n2138) );
  INVXL U2914 ( .A(n2128), .Y(n2132) );
  AOI221XL U2915 ( .A0(n2133), .A1(n2132), .B0(n2131), .B1(n2132), .C0(n2130), 
        .Y(n2136) );
  INVXL U2916 ( .A(n2134), .Y(n2135) );
  AOI221XL U2917 ( .A0(n2138), .A1(n2137), .B0(n2136), .B1(n2137), .C0(n2135), 
        .Y(n2140) );
  INVXL U2918 ( .A(n2684), .Y(n2717) );
  OAI22XL U2919 ( .A0(n2870), .A1(n2155), .B0(n2563), .B1(n2556), .Y(n1561) );
  INVXL U2920 ( .A(array_look_back[115]), .Y(n2849) );
  OAI22XL U2921 ( .A0(n2849), .A1(n2155), .B0(n2563), .B1(n2564), .Y(n1496) );
  INVXL U2922 ( .A(array_look_back[110]), .Y(n2825) );
  OAI22XL U2923 ( .A0(n2563), .A1(n2559), .B0(n2825), .B1(n2155), .Y(n1532) );
  INVXL U2924 ( .A(array_look_back[111]), .Y(n2961) );
  OAI22XL U2925 ( .A0(n2563), .A1(n2558), .B0(n2961), .B1(n2155), .Y(n1544) );
  INVXL U2926 ( .A(array_look_back[14]), .Y(n2826) );
  OAI22XL U2927 ( .A0(n2166), .A1(n2826), .B0(n2566), .B1(n2559), .Y(n1540) );
  OAI22XL U2928 ( .A0(n2166), .A1(n2869), .B0(n2566), .B1(n2556), .Y(n1593) );
  INVXL U2929 ( .A(array_look_back[19]), .Y(n2850) );
  OAI22XL U2930 ( .A0(n2166), .A1(n2850), .B0(n2566), .B1(n2564), .Y(n1504) );
  INVXL U2931 ( .A(array_look_back[139]), .Y(n2848) );
  OAI22XL U2932 ( .A0(n2848), .A1(n2164), .B0(n2171), .B1(n2564), .Y(n1494) );
  INVXL U2933 ( .A(array_look_back[143]), .Y(n2867) );
  OAI22XL U2934 ( .A0(n2867), .A1(n2164), .B0(n2171), .B1(n2556), .Y(n1681) );
  INVXL U2935 ( .A(array_look_back[140]), .Y(n2895) );
  OAI22XL U2936 ( .A0(n2895), .A1(n2164), .B0(n2171), .B1(n2554), .Y(n1556) );
  INVXL U2937 ( .A(array_look_back[116]), .Y(n2896) );
  OAI22XL U2938 ( .A0(n2896), .A1(n2155), .B0(n2563), .B1(n2554), .Y(n1564) );
  INVXL U2939 ( .A(array_look_back[104]), .Y(n2894) );
  OAI22XL U2940 ( .A0(n2160), .A1(n2894), .B0(n2580), .B1(n2554), .Y(n1568) );
  INVXL U2941 ( .A(array_look_back[138]), .Y(n2913) );
  OAI22XL U2942 ( .A0(n2913), .A1(n2164), .B0(n2171), .B1(n2567), .Y(n1482) );
  INVXL U2943 ( .A(array_look_back[114]), .Y(n2912) );
  OAI22XL U2944 ( .A0(n2912), .A1(n2155), .B0(n2563), .B1(n2567), .Y(n1484) );
  INVXL U2945 ( .A(array_look_back[117]), .Y(n2880) );
  OAI22XL U2946 ( .A0(n2880), .A1(n2155), .B0(n2563), .B1(n2555), .Y(n1563) );
  INVXL U2947 ( .A(array_look_back[141]), .Y(n2879) );
  OAI22XL U2948 ( .A0(n2879), .A1(n2164), .B0(n2171), .B1(n2555), .Y(n1555) );
  INVXL U2949 ( .A(array_look_back[21]), .Y(n2881) );
  OAI22XL U2950 ( .A0(n2166), .A1(n2881), .B0(n2566), .B1(n2555), .Y(n1595) );
  OAI22XL U2951 ( .A0(n3007), .A1(n2151), .B0(n2569), .B1(n2555), .Y(n1599) );
  INVXL U2952 ( .A(array_look_back[136]), .Y(n2933) );
  OAI22XL U2953 ( .A0(n2933), .A1(n2164), .B0(n2171), .B1(n2579), .Y(n1458) );
  INVXL U2954 ( .A(array_look_back[112]), .Y(n2934) );
  OAI22XL U2955 ( .A0(n2934), .A1(n2155), .B0(n2563), .B1(n2579), .Y(n1460) );
  INVXL U2956 ( .A(array_look_back[16]), .Y(n2935) );
  OAI22XL U2957 ( .A0(n2166), .A1(n2935), .B0(n2566), .B1(n2579), .Y(n1468) );
  INVXL U2958 ( .A(array_look_back[113]), .Y(n2923) );
  OAI22XL U2959 ( .A0(n2923), .A1(n2155), .B0(n2563), .B1(n2568), .Y(n1472) );
  INVXL U2960 ( .A(array_look_back[109]), .Y(n2945) );
  OAI22XL U2961 ( .A0(n2945), .A1(n2155), .B0(n2563), .B1(n2560), .Y(n1520) );
  INVXL U2962 ( .A(array_look_back[17]), .Y(n2924) );
  OAI22XL U2963 ( .A0(n2166), .A1(n2924), .B0(n2566), .B1(n2568), .Y(n1480) );
  INVXL U2964 ( .A(array_look_back[13]), .Y(n2947) );
  OAI22XL U2965 ( .A0(n2166), .A1(n2947), .B0(n2566), .B1(n2560), .Y(n1528) );
  INVXL U2966 ( .A(array_look_back[137]), .Y(n2921) );
  OAI22XL U2967 ( .A0(n2921), .A1(n2164), .B0(n2171), .B1(n2568), .Y(n1470) );
  INVXL U2968 ( .A(array_look_back[133]), .Y(n2944) );
  OAI22XL U2969 ( .A0(n2944), .A1(n2164), .B0(n2171), .B1(n2560), .Y(n1518) );
  INVXL U2970 ( .A(array_look_back[134]), .Y(n2824) );
  OAI22XL U2971 ( .A0(n2171), .A1(n2559), .B0(n2824), .B1(n2164), .Y(n1530) );
  INVXL U2972 ( .A(array_look_back[135]), .Y(n2959) );
  OAI22XL U2973 ( .A0(n2171), .A1(n2558), .B0(n2959), .B1(n2164), .Y(n1542) );
  INVXL U2974 ( .A(array_look_back[127]), .Y(n2847) );
  OAI22XL U2975 ( .A0(n2847), .A1(n2162), .B0(n2202), .B1(n2564), .Y(n1495) );
  INVXL U2976 ( .A(array_look_back[131]), .Y(n2868) );
  OAI22XL U2977 ( .A0(n2868), .A1(n2162), .B0(n2202), .B1(n2556), .Y(n1557) );
  INVXL U2978 ( .A(array_look_back[125]), .Y(n2922) );
  OAI22XL U2979 ( .A0(n2922), .A1(n2162), .B0(n2202), .B1(n2568), .Y(n1471) );
  INVXL U2980 ( .A(array_look_back[126]), .Y(n2910) );
  OAI22XL U2981 ( .A0(n2910), .A1(n2162), .B0(n2202), .B1(n2567), .Y(n1483) );
  INVXL U2982 ( .A(array_look_back[121]), .Y(n2943) );
  OAI22XL U2983 ( .A0(n2943), .A1(n2162), .B0(n2202), .B1(n2560), .Y(n1519) );
  INVXL U2984 ( .A(array_look_back[124]), .Y(n2932) );
  OAI22XL U2985 ( .A0(n2932), .A1(n2162), .B0(n2202), .B1(n2579), .Y(n1459) );
  INVXL U2986 ( .A(array_look_back[129]), .Y(n2878) );
  OAI22XL U2987 ( .A0(n2878), .A1(n2162), .B0(n2202), .B1(n2555), .Y(n1559) );
  INVXL U2988 ( .A(array_look_back[128]), .Y(n2893) );
  OAI22XL U2989 ( .A0(n2893), .A1(n2162), .B0(n2202), .B1(n2554), .Y(n1560) );
  INVXL U2990 ( .A(array_look_back[123]), .Y(n2957) );
  OAI22XL U2991 ( .A0(n2202), .A1(n2558), .B0(n2957), .B1(n2162), .Y(n1543) );
  INVXL U2992 ( .A(array_look_back[122]), .Y(n2823) );
  OAI22XL U2993 ( .A0(n2202), .A1(n2559), .B0(n2823), .B1(n2162), .Y(n1531) );
  INVXL U2994 ( .A(array_look_back[132]), .Y(n2976) );
  OAI22XL U2995 ( .A0(n2976), .A1(n2164), .B0(n2171), .B1(n2562), .Y(n1506) );
  INVXL U2996 ( .A(array_look_back[120]), .Y(n2972) );
  OAI22XL U2997 ( .A0(n2972), .A1(n2162), .B0(n2202), .B1(n2562), .Y(n1507) );
  INVXL U2998 ( .A(array_look_back[96]), .Y(n2974) );
  OAI22XL U2999 ( .A0(n2160), .A1(n2974), .B0(n2580), .B1(n2562), .Y(n1509) );
  INVXL U3000 ( .A(array_look_back[130]), .Y(n2163) );
  OAI22XL U3001 ( .A0(n2163), .A1(n2162), .B0(n2202), .B1(n2557), .Y(n1558) );
  INVXL U3002 ( .A(array_look_back[142]), .Y(n2165) );
  OAI22XL U3003 ( .A0(n2165), .A1(n2164), .B0(n2171), .B1(n2557), .Y(n1554) );
  INVXL U3004 ( .A(array_look_back[34]), .Y(n2859) );
  OAI22XL U3005 ( .A0(n2571), .A1(n2557), .B0(n2859), .B1(n2178), .Y(n1590) );
  INVXL U3006 ( .A(array_look_back[31]), .Y(n2844) );
  OAI22XL U3007 ( .A0(n2571), .A1(n2564), .B0(n2844), .B1(n2178), .Y(n1503) );
  INVXL U3008 ( .A(array_look_back[30]), .Y(n2908) );
  OAI22XL U3009 ( .A0(n2571), .A1(n2567), .B0(n2908), .B1(n2178), .Y(n1491) );
  INVXL U3010 ( .A(array_look_back[27]), .Y(n2956) );
  OAI22XL U3011 ( .A0(n2571), .A1(n2558), .B0(n2956), .B1(n2178), .Y(n1551) );
  NAND2XL U3012 ( .A(n2173), .B(x_array[11]), .Y(n2172) );
  OAI21XL U3013 ( .A0(n2822), .A1(n2173), .B0(n2172), .Y(n1612) );
  INVX1 U3014 ( .A(n2440), .Y(n2660) );
  NOR2X2 U3015 ( .A(n2197), .B(n2220), .Y(n2311) );
  NAND2XL U3016 ( .A(n2177), .B(x_array[2]), .Y(n2176) );
  OAI21XL U3017 ( .A0(n2822), .A1(n2177), .B0(n2176), .Y(n1603) );
  INVXL U3018 ( .A(array_look_back[39]), .Y(n2958) );
  OAI22XL U3019 ( .A0(n2573), .A1(n2558), .B0(n2958), .B1(n2423), .Y(n1550) );
  INVXL U3020 ( .A(array_look_back[44]), .Y(n2892) );
  OAI22XL U3021 ( .A0(n2573), .A1(n2554), .B0(n2892), .B1(n2423), .Y(n1588) );
  INVXL U3022 ( .A(array_look_back[36]), .Y(n2970) );
  OAI22XL U3023 ( .A0(n2573), .A1(n2562), .B0(n2970), .B1(n2423), .Y(n1514) );
  INVXL U3024 ( .A(array_look_back[42]), .Y(n2911) );
  OAI22XL U3025 ( .A0(n2573), .A1(n2567), .B0(n2911), .B1(n2423), .Y(n1490) );
  NAND2XL U3026 ( .A(n2662), .B(n2440), .Y(n2180) );
  NOR2X2 U3027 ( .A(n2180), .B(n2220), .Y(n2303) );
  NAND2XL U3028 ( .A(n2184), .B(x_array[3]), .Y(n2183) );
  OAI21XL U3029 ( .A0(n2822), .A1(n2184), .B0(n2183), .Y(n1604) );
  NAND2XL U3030 ( .A(n2187), .B(x_array[7]), .Y(n2186) );
  OAI21XL U3031 ( .A0(n2822), .A1(n2187), .B0(n2186), .Y(n1608) );
  NAND2XL U3032 ( .A(n2192), .B(n2660), .Y(n2221) );
  NOR2X1 U3033 ( .A(n2441), .B(n2221), .Y(n2312) );
  NAND2XL U3034 ( .A(n2191), .B(x_array[8]), .Y(n2190) );
  OAI21XL U3035 ( .A0(n2822), .A1(n2191), .B0(n2190), .Y(n1609) );
  NAND2XL U3036 ( .A(n2192), .B(n2440), .Y(n2212) );
  NOR2X2 U3037 ( .A(n2207), .B(n2212), .Y(n2305) );
  INVXL U3038 ( .A(n2697), .Y(n2396) );
  NAND2XL U3039 ( .A(n2196), .B(x_array[5]), .Y(n2195) );
  OAI21XL U3040 ( .A0(n2822), .A1(n2196), .B0(n2195), .Y(n1606) );
  NAND2XL U3041 ( .A(n2201), .B(x_array[6]), .Y(n2200) );
  OAI21XL U3042 ( .A0(n2822), .A1(n2201), .B0(n2200), .Y(n1607) );
  NAND2XL U3043 ( .A(n2206), .B(x_array[10]), .Y(n2205) );
  OAI21XL U3044 ( .A0(n2822), .A1(n2206), .B0(n2205), .Y(n1611) );
  NOR2X2 U3045 ( .A(n2207), .B(n2221), .Y(n2306) );
  NAND2XL U3046 ( .A(n2211), .B(x_array[4]), .Y(n2210) );
  OAI21XL U3047 ( .A0(n2822), .A1(n2211), .B0(n2210), .Y(n1605) );
  NAND2XL U3048 ( .A(n2215), .B(x_array[1]), .Y(n2214) );
  OAI21XL U3049 ( .A0(n2822), .A1(n2215), .B0(n2214), .Y(n1602) );
  NAND2XL U3050 ( .A(n2219), .B(x_array[9]), .Y(n2218) );
  OAI21XL U3051 ( .A0(n2822), .A1(n2219), .B0(n2218), .Y(n1610) );
  NOR2X2 U3052 ( .A(n2221), .B(n2220), .Y(n2314) );
  OAI211XL U3053 ( .A0(n2692), .A1(n2569), .B0(n2792), .C0(n3077), .Y(n2223)
         );
  NAND2XL U3054 ( .A(n2225), .B(x_array[0]), .Y(n2224) );
  OAI21XL U3055 ( .A0(n2822), .A1(n2225), .B0(n2224), .Y(n1601) );
  AOI22XL U3056 ( .A0(array_look_back[117]), .A1(n2308), .B0(
        array_look_back[105]), .B1(n2312), .Y(n2238) );
  AOI22XL U3057 ( .A0(array_look_back[33]), .A1(n2311), .B0(
        array_look_back[45]), .B1(n2303), .Y(n2236) );
  AOI22XL U3058 ( .A0(array_look_back[21]), .A1(n2313), .B0(
        array_look_back[141]), .B1(n2304), .Y(n2235) );
  AOI22XL U3059 ( .A0(array_look_back[69]), .A1(n2305), .B0(
        array_look_back[93]), .B1(n2309), .Y(n2234) );
  AOI22XL U3060 ( .A0(array_look_back[9]), .A1(n2314), .B0(array_look_back[57]), .B1(n2306), .Y(n2233) );
  AND4X2 U3061 ( .A(n2236), .B(n2235), .C(n2234), .D(n2233), .Y(n2237) );
  AND3X2 U3062 ( .A(n2239), .B(n2238), .C(n2237), .Y(n2334) );
  AOI22XL U3063 ( .A0(array_look_back[56]), .A1(n2306), .B0(array_look_back[8]), .B1(n2314), .Y(n2243) );
  AOI22XL U3064 ( .A0(array_look_back[68]), .A1(n2305), .B0(
        array_look_back[92]), .B1(n2309), .Y(n2241) );
  AOI22XL U3065 ( .A0(array_look_back[32]), .A1(n2311), .B0(
        array_look_back[44]), .B1(n2303), .Y(n2240) );
  AND4X2 U3066 ( .A(n2243), .B(n2242), .C(n2241), .D(n2240), .Y(n2245) );
  AOI22XL U3067 ( .A0(array_look_back[116]), .A1(n2308), .B0(
        array_look_back[104]), .B1(n2312), .Y(n2244) );
  AND3X2 U3068 ( .A(n2246), .B(n2245), .C(n2244), .Y(n2332) );
  AOI22XL U3069 ( .A0(array_look_back[46]), .A1(n2303), .B0(
        array_look_back[58]), .B1(n2306), .Y(n2249) );
  AOI22XL U3070 ( .A0(array_look_back[34]), .A1(n2311), .B0(
        array_look_back[142]), .B1(n2304), .Y(n2248) );
  AOI211X1 U3071 ( .A0(array_look_back[11]), .A1(n2314), .B0(n2260), .C0(n2259), .Y(n2325) );
  AND4X2 U3072 ( .A(n2271), .B(n2270), .C(n2269), .D(n2268), .Y(n2272) );
  INVXL U3073 ( .A(n2348), .Y(n2341) );
  INVXL U3074 ( .A(array_look_back[68]), .Y(n2890) );
  INVXL U3075 ( .A(array_look_back[69]), .Y(n2427) );
  INVXL U3076 ( .A(array_look_back[71]), .Y(n2428) );
  INVXL U3077 ( .A(array_look_back[67]), .Y(n2845) );
  INVXL U3078 ( .A(array_look_back[60]), .Y(n2429) );
  INVXL U3079 ( .A(array_look_back[70]), .Y(n2430) );
  INVXL U3080 ( .A(array_look_back[64]), .Y(n2431) );
  INVXL U3081 ( .A(array_look_back[61]), .Y(n2432) );
  INVXL U3082 ( .A(array_look_back[63]), .Y(n2433) );
  INVXL U3083 ( .A(array_look_back[66]), .Y(n2434) );
  INVXL U3084 ( .A(array_look_back[62]), .Y(n2435) );
  INVXL U3085 ( .A(array_look_back[65]), .Y(n2437) );
  INVXL U3086 ( .A(array_look_back[80]), .Y(n2891) );
  INVXL U3087 ( .A(array_look_back[82]), .Y(n2858) );
  INVXL U3088 ( .A(array_look_back[79]), .Y(n2843) );
  INVXL U3089 ( .A(array_look_back[78]), .Y(n2909) );
  INVXL U3090 ( .A(array_look_back[75]), .Y(n2955) );
  AOI222XL U3091 ( .A0(n2683), .A1(n2467), .B0(n2683), .B1(n2464), .C0(n2467), 
        .C1(n2464), .Y(n2492) );
  INVXL U3092 ( .A(array_look_back[88]), .Y(n2500) );
  INVXL U3093 ( .A(array_look_back[94]), .Y(n2501) );
  INVXL U3094 ( .A(array_look_back[89]), .Y(n2502) );
  INVXL U3095 ( .A(array_look_back[93]), .Y(n2503) );
  INVXL U3096 ( .A(array_look_back[85]), .Y(n2504) );
  INVXL U3097 ( .A(array_look_back[91]), .Y(n2846) );
  INVXL U3098 ( .A(array_look_back[92]), .Y(n2899) );
  INVXL U3099 ( .A(array_look_back[90]), .Y(n2505) );
  INVXL U3100 ( .A(array_look_back[95]), .Y(n2506) );
  INVXL U3101 ( .A(array_look_back[86]), .Y(n2513) );
  INVXL U3102 ( .A(array_look_back[84]), .Y(n2514) );
  INVXL U3103 ( .A(array_look_back[87]), .Y(n2516) );
  INVXL U3104 ( .A(count_out[2]), .Y(n2835) );
  AOI221XL U3105 ( .A0(count_out[2]), .A1(n2832), .B0(n2835), .B1(n2526), .C0(
        n3086), .Y(N6084) );
  OAI2BB2XL U3106 ( .B0(n2529), .B1(n3086), .A0N(n2528), .A1N(n2527), .Y(n1683) );
  AOI2BB1XL U3107 ( .A0N(in_valid), .A1N(count_receive[0]), .B0(n2530), .Y(
        n1679) );
  OAI2BB2XL U3108 ( .B0(n3007), .B1(n2533), .A0N(n2532), .A1N(n2531), .Y(n1675) );
  OAI2BB2XL U3109 ( .B0(n2537), .B1(n2534), .A0N(n2792), .A1N(array_in[1]), 
        .Y(n1674) );
  NAND2XL U3110 ( .A(col[1]), .B(col[3]), .Y(n2536) );
  OAI2BB2XL U3111 ( .B0(n2537), .B1(n2536), .A0N(n2792), .A1N(array_in[11]), 
        .Y(n1664) );
  OAI2BB1XL U3112 ( .A0N(count[3]), .A1N(n2538), .B0(n2792), .Y(n1662) );
  OAI2BB2XL U3113 ( .B0(n2569), .B1(n2554), .A0N(n2792), .A1N(
        array_look_back[8]), .Y(n1600) );
  OAI2BB2XL U3114 ( .B0(n2569), .B1(n2557), .A0N(n2792), .A1N(
        array_look_back[10]), .Y(n1598) );
  OAI2BB2XL U3115 ( .B0(n2566), .B1(n2554), .A0N(n2565), .A1N(
        array_look_back[20]), .Y(n1596) );
  OAI2BB2XL U3116 ( .B0(n2566), .B1(n2557), .A0N(n2565), .A1N(
        array_look_back[22]), .Y(n1594) );
  OAI2BB2XL U3117 ( .B0(n2580), .B1(n2555), .A0N(n2578), .A1N(
        array_look_back[105]), .Y(n1567) );
  OAI2BB2XL U3118 ( .B0(n2580), .B1(n2557), .A0N(n2578), .A1N(
        array_look_back[106]), .Y(n1566) );
  OAI2BB2XL U3119 ( .B0(n2563), .B1(n2557), .A0N(array_look_back[118]), .A1N(
        n2561), .Y(n1562) );
  OAI2BB2XL U3120 ( .B0(n2569), .B1(n2558), .A0N(n2792), .A1N(
        array_look_back[3]), .Y(n1553) );
  OAI2BB2XL U3121 ( .B0(n2566), .B1(n2558), .A0N(n2565), .A1N(
        array_look_back[15]), .Y(n1552) );
  OAI2BB2XL U3122 ( .B0(n2580), .B1(n2558), .A0N(n2578), .A1N(
        array_look_back[99]), .Y(n1545) );
  OAI2BB2XL U3123 ( .B0(n2569), .B1(n2559), .A0N(n2792), .A1N(
        array_look_back[2]), .Y(n1541) );
  OAI2BB2XL U3124 ( .B0(n2571), .B1(n2559), .A0N(array_look_back[26]), .A1N(
        n2570), .Y(n1539) );
  OAI2BB2XL U3125 ( .B0(n2580), .B1(n2559), .A0N(n2578), .A1N(
        array_look_back[98]), .Y(n1533) );
  OAI2BB2XL U3126 ( .B0(n2569), .B1(n2560), .A0N(n2792), .A1N(
        array_look_back[1]), .Y(n1529) );
  OAI2BB2XL U3127 ( .B0(n2580), .B1(n2560), .A0N(n2578), .A1N(
        array_look_back[97]), .Y(n1521) );
  OAI2BB2XL U3128 ( .B0(n2569), .B1(n2562), .A0N(n2792), .A1N(
        array_look_back[0]), .Y(n1517) );
  OAI2BB2XL U3129 ( .B0(n2566), .B1(n2562), .A0N(n2565), .A1N(
        array_look_back[12]), .Y(n1516) );
  OAI2BB2XL U3130 ( .B0(n2571), .B1(n2562), .A0N(array_look_back[24]), .A1N(
        n2570), .Y(n1515) );
  OAI2BB2XL U3131 ( .B0(n2563), .B1(n2562), .A0N(array_look_back[108]), .A1N(
        n2561), .Y(n1508) );
  OAI2BB2XL U3132 ( .B0(n2569), .B1(n2564), .A0N(n2792), .A1N(
        array_look_back[7]), .Y(n1505) );
  OAI2BB2XL U3133 ( .B0(n2580), .B1(n2564), .A0N(n2578), .A1N(
        array_look_back[103]), .Y(n1497) );
  OAI2BB2XL U3134 ( .B0(n2569), .B1(n2568), .A0N(n2792), .A1N(
        array_look_back[5]), .Y(n1481) );
  OAI2BB2XL U3135 ( .B0(n2580), .B1(n2568), .A0N(n2578), .A1N(
        array_look_back[101]), .Y(n1473) );
  OAI2BB2XL U3136 ( .B0(n2569), .B1(n2579), .A0N(n2792), .A1N(
        array_look_back[4]), .Y(n1469) );
  OAI2BB2XL U3137 ( .B0(n2580), .B1(n2579), .A0N(n2578), .A1N(
        array_look_back[100]), .Y(n1461) );
  INVXL U3138 ( .A(sub_array[11]), .Y(n2588) );
  INVXL U3139 ( .A(sub_array[12]), .Y(n2590) );
  INVXL U3140 ( .A(sub_array[14]), .Y(n2601) );
  INVXL U3141 ( .A(sub_array[15]), .Y(n2615) );
  INVXL U3142 ( .A(sub_array[18]), .Y(n2627) );
  INVXL U3143 ( .A(sub_array[21]), .Y(n2637) );
  INVXL U3144 ( .A(sub_array[5]), .Y(n2643) );
  INVXL U3145 ( .A(sub_array[9]), .Y(n2658) );
  AOI222X1 U3146 ( .A0(n2671), .A1(n2662), .B0(n2671), .B1(n2661), .C0(n2662), 
        .C1(n2661), .Y(n2668) );
  AOI222X1 U3147 ( .A0(n2207), .A1(n2663), .B0(n2207), .B1(n2668), .C0(n2663), 
        .C1(n2668), .Y(n2665) );
  XOR2X1 U3148 ( .A(n2665), .B(n2664), .Y(n2745) );
  AOI222X1 U3149 ( .A0(n2665), .A1(n2667), .B0(n2665), .B1(n2666), .C0(n2667), 
        .C1(n2666), .Y(n2759) );
  AOI222XL U3150 ( .A0(n2683), .A1(x[2]), .B0(n2683), .B1(n2689), .C0(x[2]), 
        .C1(n2689), .Y(n2715) );
  AOI222XL U3151 ( .A0(n2708), .A1(n2801), .B0(n2800), .B1(n2707), .C0(n2706), 
        .C1(n2799), .Y(n2691) );
  NAND2XL U3152 ( .A(n2691), .B(add_array[0]), .Y(n2690) );
  OAI21XL U3153 ( .A0(n2822), .A1(n2691), .B0(n2690), .Y(n1430) );
  INVXL U3154 ( .A(add_array[2]), .Y(n2694) );
  AOI222XL U3155 ( .A0(n2708), .A1(n2806), .B0(n2707), .B1(n2805), .C0(n2804), 
        .C1(n2706), .Y(n2693) );
  AOI222XL U3156 ( .A0(n2708), .A1(n2811), .B0(n2707), .B1(n2810), .C0(n2809), 
        .C1(n2706), .Y(n2701) );
  NAND2XL U3157 ( .A(n2701), .B(add_array[4]), .Y(n2700) );
  OAI21XL U3158 ( .A0(n2822), .A1(n2701), .B0(n2700), .Y(n1428) );
  INVX1 U3159 ( .A(n2759), .Y(n2794) );
  INVXL U3160 ( .A(n2744), .Y(n2730) );
  OAI31XL U3161 ( .A0(n2794), .A1(n2745), .A2(n2730), .B0(n2792), .Y(n2727) );
  AOI222XL U3162 ( .A0(n2713), .A1(n2711), .B0(n2713), .B1(n3081), .C0(n2711), 
        .C1(n3081), .Y(n2767) );
  XOR2XL U3163 ( .A(n2714), .B(n2715), .Y(n2763) );
  INVXL U3164 ( .A(n2715), .Y(n2716) );
  AOI222XL U3165 ( .A0(N4586), .A1(n2717), .B0(N4586), .B1(n2716), .C0(n2717), 
        .C1(n2716), .Y(n2762) );
  AOI222XL U3166 ( .A0(n2727), .A1(n2801), .B0(n2800), .B1(n2726), .C0(n2799), 
        .C1(n2725), .Y(n2719) );
  INVXL U3167 ( .A(add_array[10]), .Y(n2722) );
  AOI222XL U3168 ( .A0(n2727), .A1(n2806), .B0(n2805), .B1(n2726), .C0(n2804), 
        .C1(n2725), .Y(n2721) );
  AOI222XL U3169 ( .A0(n2727), .A1(n2811), .B0(n2810), .B1(n2726), .C0(n2809), 
        .C1(n2725), .Y(n2723) );
  INVXL U3170 ( .A(add_array[14]), .Y(n2729) );
  AOI222XL U3171 ( .A0(n2727), .A1(n2818), .B0(n2817), .B1(n2726), .C0(n2725), 
        .C1(n2814), .Y(n2728) );
  NAND2XL U3172 ( .A(n2745), .B(n2730), .Y(n2761) );
  OAI21XL U3173 ( .A0(n2794), .A1(n2761), .B0(n2792), .Y(n2741) );
  AOI222XL U3174 ( .A0(n2741), .A1(n2801), .B0(n2800), .B1(n2740), .C0(n2799), 
        .C1(n2739), .Y(n2734) );
  NAND2XL U3175 ( .A(n2734), .B(add_array[1]), .Y(n2733) );
  OAI21XL U3176 ( .A0(n2822), .A1(n2734), .B0(n2733), .Y(n1422) );
  AOI222XL U3177 ( .A0(n2741), .A1(n2806), .B0(n2805), .B1(n2740), .C0(n2804), 
        .C1(n2739), .Y(n2736) );
  NAND2XL U3178 ( .A(n2736), .B(add_array[3]), .Y(n2735) );
  OAI21XL U3179 ( .A0(n2822), .A1(n2736), .B0(n2735), .Y(n1421) );
  AOI222XL U3180 ( .A0(n2741), .A1(n2811), .B0(n2810), .B1(n2740), .C0(n2809), 
        .C1(n2739), .Y(n2737) );
  INVXL U3181 ( .A(add_array[7]), .Y(n2743) );
  AOI222XL U3182 ( .A0(n2741), .A1(n2818), .B0(n2817), .B1(n2740), .C0(n2739), 
        .C1(n2814), .Y(n2742) );
  INVXL U3183 ( .A(add_array[9]), .Y(n2749) );
  OAI31XL U3184 ( .A0(n2794), .A1(n2745), .A2(n2744), .B0(n2792), .Y(n2756) );
  AOI222XL U3185 ( .A0(n2756), .A1(n2801), .B0(n2800), .B1(n2755), .C0(n2799), 
        .C1(n2754), .Y(n2748) );
  INVXL U3186 ( .A(add_array[11]), .Y(n2751) );
  AOI222XL U3187 ( .A0(n2756), .A1(n2806), .B0(n2805), .B1(n2755), .C0(n2804), 
        .C1(n2754), .Y(n2750) );
  AOI222XL U3188 ( .A0(n2756), .A1(n2811), .B0(n2810), .B1(n2755), .C0(n2809), 
        .C1(n2754), .Y(n2752) );
  INVXL U3189 ( .A(add_array[15]), .Y(n2758) );
  AOI222XL U3190 ( .A0(n2756), .A1(n2818), .B0(n2817), .B1(n2755), .C0(n2754), 
        .C1(n2814), .Y(n2757) );
  OAI31XL U3191 ( .A0(n2761), .A1(n2760), .A2(n2759), .B0(n2792), .Y(n2784) );
  AOI222XL U3192 ( .A0(n2771), .A1(n2784), .B0(n2770), .B1(n2782), .C0(n2769), 
        .C1(n2787), .Y(n2772) );
  INVXL U3193 ( .A(add_array[19]), .Y(n2780) );
  AOI22XL U3194 ( .A0(n2784), .A1(n2775), .B0(n2787), .B1(n2774), .Y(n2776) );
  OAI21XL U3195 ( .A0(n2778), .A1(n2777), .B0(n2776), .Y(n2779) );
  AOI22XL U3196 ( .A0(n2784), .A1(n2783), .B0(n2782), .B1(n2781), .Y(n2785) );
  AOI31XL U3197 ( .A0(n2789), .A1(n2788), .A2(n2787), .B0(n2786), .Y(n2790) );
  AOI222XL U3198 ( .A0(n2819), .A1(n2801), .B0(n2800), .B1(n2816), .C0(n2799), 
        .C1(n2815), .Y(n2802) );
  INVXL U3199 ( .A(add_array[18]), .Y(n2808) );
  AOI222XL U3200 ( .A0(n2819), .A1(n2806), .B0(n2805), .B1(n2816), .C0(n2804), 
        .C1(n2815), .Y(n2807) );
  AOI222XL U3201 ( .A0(n2819), .A1(n2811), .B0(n2810), .B1(n2816), .C0(n2809), 
        .C1(n2815), .Y(n2813) );
  NAND2XL U3202 ( .A(n2813), .B(add_array[20]), .Y(n2812) );
  OAI21XL U3203 ( .A0(n2822), .A1(n2813), .B0(n2812), .Y(n1409) );
  AOI222XL U3204 ( .A0(n2819), .A1(n2818), .B0(n2817), .B1(n2816), .C0(n2815), 
        .C1(n2814), .Y(n2821) );
  NAND2XL U3205 ( .A(n2821), .B(add_array[22]), .Y(n2820) );
  OAI21XL U3206 ( .A0(n2822), .A1(n2821), .B0(n2820), .Y(n1408) );
  NAND2XL U3207 ( .A(count_out[3]), .B(n3085), .Y(n2831) );
  INVXL U3208 ( .A(n3052), .Y(n2971) );
  OAI22XL U3209 ( .A0(n2824), .A1(n2975), .B0(n2823), .B1(n2971), .Y(n2842) );
  NAND2XL U3210 ( .A(count_out[0]), .B(n2830), .Y(n2829) );
  INVXL U3211 ( .A(n3058), .Y(n2946) );
  NAND3XL U3212 ( .A(n2827), .B(count_out[0]), .C(count_out[3]), .Y(n2960) );
  OAI22XL U3213 ( .A0(n2826), .A1(n2946), .B0(n2825), .B1(n2960), .Y(n2841) );
  NOR3XL U3214 ( .A(count_out[0]), .B(count_out[3]), .C(n2827), .Y(n2828) );
  NAND2XL U3215 ( .A(n2828), .B(n2835), .Y(n2984) );
  INVXL U3216 ( .A(n2984), .Y(n3062) );
  NAND2XL U3217 ( .A(count_out[2]), .B(n2828), .Y(n2986) );
  INVXL U3218 ( .A(n2986), .Y(n3060) );
  AOI22XL U3219 ( .A0(array_look_back[26]), .A1(n3062), .B0(
        array_look_back[74]), .B1(n3060), .Y(n2839) );
  AOI22XL U3220 ( .A0(array_look_back[86]), .A1(n3059), .B0(
        array_look_back[62]), .B1(n3061), .Y(n2838) );
  NAND2XL U3221 ( .A(n2830), .B(n3085), .Y(n2834) );
  AOI22XL U3222 ( .A0(array_look_back[2]), .A1(n3053), .B0(array_look_back[98]), .B1(n3055), .Y(n2837) );
  NAND3XL U3223 ( .A(n2835), .B(n2833), .C(n2832), .Y(n2969) );
  INVXL U3224 ( .A(n2969), .Y(n3054) );
  AOI22XL U3225 ( .A0(array_look_back[38]), .A1(n3054), .B0(
        array_look_back[50]), .B1(n3051), .Y(n2836) );
  NAND4XL U3226 ( .A(n2839), .B(n2838), .C(n2837), .D(n2836), .Y(n2840) );
  NOR3XL U3227 ( .A(n2842), .B(n2841), .C(n2840), .Y(n3032) );
  AOI22XL U3228 ( .A0(array_look_back[7]), .A1(n3053), .B0(
        array_look_back[103]), .B1(n3055), .Y(n2857) );
  AOI22XL U3229 ( .A0(array_look_back[43]), .A1(n3054), .B0(
        array_look_back[55]), .B1(n3051), .Y(n2856) );
  OAI22XL U3230 ( .A0(n2844), .A1(n2984), .B0(n2843), .B1(n2986), .Y(n2854) );
  INVXL U3231 ( .A(n3061), .Y(n2889) );
  OAI22XL U3232 ( .A0(n2846), .A1(n2898), .B0(n2845), .B1(n2889), .Y(n2853) );
  OAI22XL U3233 ( .A0(n2848), .A1(n2975), .B0(n2847), .B1(n2971), .Y(n2852) );
  OAI22XL U3234 ( .A0(n2850), .A1(n2946), .B0(n2849), .B1(n2960), .Y(n2851) );
  NOR4XL U3235 ( .A(n2854), .B(n2853), .C(n2852), .D(n2851), .Y(n2855) );
  NAND3XL U3236 ( .A(n2857), .B(n2856), .C(n2855), .Y(n3010) );
  AOI22XL U3237 ( .A0(array_look_back[94]), .A1(n3059), .B0(
        array_look_back[70]), .B1(n3061), .Y(n2866) );
  INVXL U3238 ( .A(n2960), .Y(n3057) );
  AOI22XL U3239 ( .A0(array_look_back[22]), .A1(n3058), .B0(
        array_look_back[118]), .B1(n3057), .Y(n2865) );
  AOI22XL U3240 ( .A0(array_look_back[10]), .A1(n3053), .B0(
        array_look_back[58]), .B1(n3051), .Y(n2864) );
  OAI22XL U3241 ( .A0(n2859), .A1(n2984), .B0(n2858), .B1(n2986), .Y(n2862) );
  AOI22XL U3242 ( .A0(array_look_back[130]), .A1(n3052), .B0(
        array_look_back[106]), .B1(n3055), .Y(n2860) );
  OAI2BB1XL U3243 ( .A0N(array_look_back[142]), .A1N(n3056), .B0(n2860), .Y(
        n2861) );
  AOI211XL U3244 ( .A0(array_look_back[46]), .A1(n3054), .B0(n2862), .C0(n2861), .Y(n2863) );
  NAND4XL U3245 ( .A(n2866), .B(n2865), .C(n2864), .D(n2863), .Y(n3049) );
  OAI22XL U3246 ( .A0(n2868), .A1(n2971), .B0(n2867), .B1(n2975), .Y(n2877) );
  OAI22XL U3247 ( .A0(n2870), .A1(n2960), .B0(n2869), .B1(n2946), .Y(n2876) );
  AOI22XL U3248 ( .A0(array_look_back[35]), .A1(n3062), .B0(
        array_look_back[83]), .B1(n3060), .Y(n2874) );
  AOI22XL U3249 ( .A0(array_look_back[95]), .A1(n3059), .B0(
        array_look_back[71]), .B1(n3061), .Y(n2873) );
  AOI22XL U3250 ( .A0(array_look_back[107]), .A1(n3055), .B0(
        array_look_back[11]), .B1(n3053), .Y(n2872) );
  AOI22XL U3251 ( .A0(array_look_back[47]), .A1(n3054), .B0(
        array_look_back[59]), .B1(n3051), .Y(n2871) );
  NAND4XL U3252 ( .A(n2874), .B(n2873), .C(n2872), .D(n2871), .Y(n2875) );
  NOR3XL U3253 ( .A(n2877), .B(n2876), .C(n2875), .Y(n3025) );
  OAI22XL U3254 ( .A0(n2879), .A1(n2975), .B0(n2878), .B1(n2971), .Y(n2888) );
  OAI22XL U3255 ( .A0(n2881), .A1(n2946), .B0(n2880), .B1(n2960), .Y(n2887) );
  AOI22XL U3256 ( .A0(array_look_back[33]), .A1(n3062), .B0(
        array_look_back[81]), .B1(n3060), .Y(n2885) );
  AOI22XL U3257 ( .A0(array_look_back[69]), .A1(n3061), .B0(
        array_look_back[93]), .B1(n3059), .Y(n2884) );
  AOI22XL U3258 ( .A0(array_look_back[9]), .A1(n3053), .B0(
        array_look_back[105]), .B1(n3055), .Y(n2883) );
  AOI22XL U3259 ( .A0(array_look_back[45]), .A1(n3054), .B0(
        array_look_back[57]), .B1(n3051), .Y(n2882) );
  NAND4XL U3260 ( .A(n2885), .B(n2884), .C(n2883), .D(n2882), .Y(n2886) );
  NOR3XL U3261 ( .A(n2888), .B(n2887), .C(n2886), .Y(n3050) );
  OAI22XL U3262 ( .A0(n2891), .A1(n2986), .B0(n2890), .B1(n2889), .Y(n2906) );
  OAI22XL U3263 ( .A0(n2893), .A1(n2971), .B0(n2892), .B1(n2969), .Y(n2905) );
  INVXL U3264 ( .A(n3055), .Y(n2973) );
  OAI22XL U3265 ( .A0(n2895), .A1(n2975), .B0(n2894), .B1(n2973), .Y(n2904) );
  INVXL U3266 ( .A(n3051), .Y(n2989) );
  AOI22XL U3267 ( .A0(array_look_back[32]), .A1(n3062), .B0(
        array_look_back[20]), .B1(n3058), .Y(n2901) );
  OAI2BB2XL U3268 ( .B0(n2896), .B1(n2960), .A0N(array_look_back[8]), .A1N(
        n3053), .Y(n2897) );
  AOI2BB1XL U3269 ( .A0N(n2899), .A1N(n2898), .B0(n2897), .Y(n2900) );
  OAI211XL U3270 ( .A0(n2902), .A1(n2989), .B0(n2901), .C0(n2900), .Y(n2903)
         );
  NOR4XL U3271 ( .A(n2906), .B(n2905), .C(n2904), .D(n2903), .Y(n2907) );
  NAND4BXL U3272 ( .AN(n3049), .B(n3025), .C(n3050), .D(n2907), .Y(n2998) );
  AOI22XL U3273 ( .A0(array_look_back[90]), .A1(n3059), .B0(
        array_look_back[66]), .B1(n3061), .Y(n2920) );
  AOI22XL U3274 ( .A0(array_look_back[102]), .A1(n3055), .B0(
        array_look_back[18]), .B1(n3058), .Y(n2919) );
  AOI22XL U3275 ( .A0(array_look_back[6]), .A1(n3053), .B0(array_look_back[54]), .B1(n3051), .Y(n2918) );
  OAI22XL U3276 ( .A0(n2909), .A1(n2986), .B0(n2908), .B1(n2984), .Y(n2916) );
  OAI22XL U3277 ( .A0(n2911), .A1(n2969), .B0(n2910), .B1(n2971), .Y(n2915) );
  OAI22XL U3278 ( .A0(n2913), .A1(n2975), .B0(n2912), .B1(n2960), .Y(n2914) );
  NOR3XL U3279 ( .A(n2916), .B(n2915), .C(n2914), .Y(n2917) );
  NAND4XL U3280 ( .A(n2920), .B(n2919), .C(n2918), .D(n2917), .Y(n3011) );
  NOR3XL U3281 ( .A(n3010), .B(n2998), .C(n3011), .Y(n3013) );
  OAI22XL U3282 ( .A0(n2922), .A1(n2971), .B0(n2921), .B1(n2975), .Y(n2931) );
  OAI22XL U3283 ( .A0(n2924), .A1(n2946), .B0(n2923), .B1(n2960), .Y(n2930) );
  AOI22XL U3284 ( .A0(array_look_back[29]), .A1(n3062), .B0(
        array_look_back[77]), .B1(n3060), .Y(n2928) );
  AOI22XL U3285 ( .A0(array_look_back[89]), .A1(n3059), .B0(
        array_look_back[65]), .B1(n3061), .Y(n2927) );
  AOI22XL U3286 ( .A0(array_look_back[5]), .A1(n3053), .B0(
        array_look_back[101]), .B1(n3055), .Y(n2926) );
  AOI22XL U3287 ( .A0(array_look_back[41]), .A1(n3054), .B0(
        array_look_back[53]), .B1(n3051), .Y(n2925) );
  NAND4XL U3288 ( .A(n2928), .B(n2927), .C(n2926), .D(n2925), .Y(n2929) );
  NOR3XL U3289 ( .A(n2931), .B(n2930), .C(n2929), .Y(n3044) );
  OAI22XL U3290 ( .A0(n2933), .A1(n2975), .B0(n2932), .B1(n2971), .Y(n2942) );
  OAI22XL U3291 ( .A0(n2935), .A1(n2946), .B0(n2934), .B1(n2960), .Y(n2941) );
  AOI22XL U3292 ( .A0(array_look_back[28]), .A1(n3062), .B0(
        array_look_back[76]), .B1(n3060), .Y(n2939) );
  AOI22XL U3293 ( .A0(array_look_back[64]), .A1(n3061), .B0(
        array_look_back[88]), .B1(n3059), .Y(n2938) );
  AOI22XL U3294 ( .A0(array_look_back[100]), .A1(n3055), .B0(
        array_look_back[4]), .B1(n3053), .Y(n2937) );
  AOI22XL U3295 ( .A0(array_look_back[52]), .A1(n3051), .B0(
        array_look_back[40]), .B1(n3054), .Y(n2936) );
  NAND4XL U3296 ( .A(n2939), .B(n2938), .C(n2937), .D(n2936), .Y(n2940) );
  NOR3XL U3297 ( .A(n2942), .B(n2941), .C(n2940), .Y(n3014) );
  NAND3XL U3298 ( .A(n3013), .B(n3044), .C(n3014), .Y(n3031) );
  INVXL U3299 ( .A(n3031), .Y(n3029) );
  AND2XL U3300 ( .A(n3032), .B(n3029), .Y(n3045) );
  OAI22XL U3301 ( .A0(n2944), .A1(n2975), .B0(n2943), .B1(n2971), .Y(n2954) );
  OAI22XL U3302 ( .A0(n2947), .A1(n2946), .B0(n2945), .B1(n2960), .Y(n2953) );
  AOI22XL U3303 ( .A0(array_look_back[25]), .A1(n3062), .B0(
        array_look_back[73]), .B1(n3060), .Y(n2951) );
  AOI22XL U3304 ( .A0(array_look_back[61]), .A1(n3061), .B0(
        array_look_back[85]), .B1(n3059), .Y(n2950) );
  AOI22XL U3305 ( .A0(array_look_back[1]), .A1(n3053), .B0(array_look_back[97]), .B1(n3055), .Y(n2949) );
  AOI22XL U3306 ( .A0(array_look_back[37]), .A1(n3054), .B0(
        array_look_back[49]), .B1(n3051), .Y(n2948) );
  NAND4XL U3307 ( .A(n2951), .B(n2950), .C(n2949), .D(n2948), .Y(n2952) );
  NOR3XL U3308 ( .A(n2954), .B(n2953), .C(n2952), .Y(n3046) );
  AOI22XL U3309 ( .A0(array_look_back[63]), .A1(n3061), .B0(
        array_look_back[87]), .B1(n3059), .Y(n2968) );
  AOI22XL U3310 ( .A0(array_look_back[99]), .A1(n3055), .B0(
        array_look_back[15]), .B1(n3058), .Y(n2967) );
  AOI22XL U3311 ( .A0(array_look_back[3]), .A1(n3053), .B0(array_look_back[51]), .B1(n3051), .Y(n2966) );
  OAI22XL U3312 ( .A0(n2956), .A1(n2984), .B0(n2955), .B1(n2986), .Y(n2964) );
  OAI22XL U3313 ( .A0(n2958), .A1(n2969), .B0(n2957), .B1(n2971), .Y(n2963) );
  OAI22XL U3314 ( .A0(n2961), .A1(n2960), .B0(n2959), .B1(n2975), .Y(n2962) );
  NOR3XL U3315 ( .A(n2964), .B(n2963), .C(n2962), .Y(n2965) );
  NAND4XL U3316 ( .A(n2968), .B(n2967), .C(n2966), .D(n2965), .Y(n3028) );
  OAI22XL U3317 ( .A0(n2972), .A1(n2971), .B0(n2970), .B1(n2969), .Y(n2983) );
  OAI22XL U3318 ( .A0(n2976), .A1(n2975), .B0(n2974), .B1(n2973), .Y(n2982) );
  AOI22XL U3319 ( .A0(array_look_back[24]), .A1(n3062), .B0(
        array_look_back[12]), .B1(n3058), .Y(n2980) );
  AOI22XL U3320 ( .A0(array_look_back[72]), .A1(n3060), .B0(
        array_look_back[60]), .B1(n3061), .Y(n2979) );
  AOI22XL U3321 ( .A0(array_look_back[48]), .A1(n3051), .B0(
        array_look_back[108]), .B1(n3057), .Y(n2978) );
  AOI22XL U3322 ( .A0(array_look_back[0]), .A1(n3053), .B0(array_look_back[84]), .B1(n3059), .Y(n2977) );
  NAND4XL U3323 ( .A(n2980), .B(n2979), .C(n2978), .D(n2977), .Y(n2981) );
  NOR4XL U3324 ( .A(n3028), .B(n2983), .C(n2982), .D(n2981), .Y(n2997) );
  AOI22XL U3325 ( .A0(array_in[5]), .A1(n3061), .B0(array_in[7]), .B1(n3059), 
        .Y(n2996) );
  AOI22XL U3326 ( .A0(array_in[10]), .A1(n3052), .B0(array_in[3]), .B1(n3054), 
        .Y(n2995) );
  AOI22XL U3327 ( .A0(array_in[9]), .A1(n3057), .B0(array_in[11]), .B1(n3056), 
        .Y(n2994) );
  OAI22XL U3328 ( .A0(n2987), .A1(n2986), .B0(n2985), .B1(n2984), .Y(n2992) );
  AOI22XL U3329 ( .A0(array_in[1]), .A1(n3058), .B0(array_in[0]), .B1(n3053), 
        .Y(n2988) );
  OAI21XL U3330 ( .A0(n2990), .A1(n2989), .B0(n2988), .Y(n2991) );
  AOI211XL U3331 ( .A0(array_in[8]), .A1(n3055), .B0(n2992), .C0(n2991), .Y(
        n2993) );
  NAND4XL U3332 ( .A(n2996), .B(n2995), .C(n2994), .D(n2993), .Y(n3067) );
  AOI31XL U3333 ( .A0(n3045), .A1(n3046), .A2(n2997), .B0(n3067), .Y(n3009) );
  INVXL U3334 ( .A(n2998), .Y(n3012) );
  AOI22XL U3335 ( .A0(n3055), .A1(row_store[35]), .B0(n3054), .B1(
        row_store[15]), .Y(n3005) );
  AOI22XL U3336 ( .A0(n3051), .A1(row_store[19]), .B0(n3053), .B1(row_store[3]), .Y(n3004) );
  AOI22XL U3337 ( .A0(n3056), .A1(row_store[47]), .B0(n3052), .B1(
        row_store[43]), .Y(n3002) );
  AOI22XL U3338 ( .A0(n3058), .A1(row_store[7]), .B0(n3057), .B1(row_store[39]), .Y(n3001) );
  AOI22XL U3339 ( .A0(n3059), .A1(row_store[31]), .B0(n3061), .B1(
        row_store[23]), .Y(n3000) );
  AOI22XL U3340 ( .A0(n3060), .A1(row_store[27]), .B0(n3062), .B1(
        row_store[11]), .Y(n2999) );
  NAND4XL U3341 ( .A(n3005), .B(n3004), .C(n3003), .D(n3067), .Y(n3006) );
  OAI2BB1XL U3342 ( .A0N(n3009), .A1N(n3012), .B0(n3006), .Y(n3008) );
  INVXL U3343 ( .A(n3086), .Y(n3072) );
  OAI2BB2XL U3344 ( .B0(n3086), .B1(n3008), .A0N(n3076), .A1N(out[3]), .Y(
        n1399) );
  OAI2BB1XL U3345 ( .A0N(n3010), .A1N(n3012), .B0(n3009), .Y(n3026) );
  NAND2XL U3346 ( .A(n3012), .B(n3011), .Y(n3030) );
  INVXL U3347 ( .A(n3013), .Y(n3043) );
  AOI32XL U3348 ( .A0(n3044), .A1(n3030), .A2(n3014), .B0(n3043), .B1(n3030), 
        .Y(n3023) );
  AOI22XL U3349 ( .A0(n3055), .A1(row_store[34]), .B0(n3054), .B1(
        row_store[14]), .Y(n3021) );
  AOI22XL U3350 ( .A0(n3051), .A1(row_store[18]), .B0(n3053), .B1(row_store[2]), .Y(n3020) );
  AOI22XL U3351 ( .A0(n3056), .A1(row_store[46]), .B0(n3052), .B1(
        row_store[42]), .Y(n3018) );
  AOI22XL U3352 ( .A0(n3058), .A1(row_store[6]), .B0(n3057), .B1(row_store[38]), .Y(n3017) );
  AOI22XL U3353 ( .A0(n3059), .A1(row_store[30]), .B0(n3061), .B1(
        row_store[22]), .Y(n3016) );
  AOI22XL U3354 ( .A0(n3060), .A1(row_store[26]), .B0(n3062), .B1(
        row_store[10]), .Y(n3015) );
  NAND4XL U3355 ( .A(n3021), .B(n3020), .C(n3019), .D(n3067), .Y(n3022) );
  OAI211XL U3356 ( .A0(n3026), .A1(n3023), .B0(n3072), .C0(n3022), .Y(n3024)
         );
  OAI2BB1XL U3357 ( .A0N(n3076), .A1N(out[2]), .B0(n3024), .Y(n1398) );
  INVXL U3358 ( .A(n3025), .Y(n3027) );
  AOI211XL U3359 ( .A0(n3029), .A1(n3028), .B0(n3027), .C0(n3026), .Y(n3048)
         );
  OAI211XL U3360 ( .A0(n3032), .A1(n3031), .B0(n3048), .C0(n3030), .Y(n3041)
         );
  AOI22XL U3361 ( .A0(n3055), .A1(row_store[33]), .B0(n3054), .B1(
        row_store[13]), .Y(n3039) );
  AOI22XL U3362 ( .A0(n3051), .A1(row_store[17]), .B0(n3053), .B1(row_store[1]), .Y(n3038) );
  AOI22XL U3363 ( .A0(n3056), .A1(row_store[45]), .B0(n3052), .B1(
        row_store[41]), .Y(n3036) );
  AOI22XL U3364 ( .A0(n3058), .A1(row_store[5]), .B0(n3057), .B1(row_store[37]), .Y(n3035) );
  AOI22XL U3365 ( .A0(n3059), .A1(row_store[29]), .B0(n3061), .B1(
        row_store[21]), .Y(n3034) );
  AOI22XL U3366 ( .A0(n3060), .A1(row_store[25]), .B0(n3062), .B1(row_store[9]), .Y(n3033) );
  NAND4XL U3367 ( .A(n3039), .B(n3038), .C(n3037), .D(n3067), .Y(n3040) );
  OAI211XL U3368 ( .A0(n3049), .A1(n3041), .B0(n3072), .C0(n3040), .Y(n3042)
         );
  OAI2BB1XL U3369 ( .A0N(n3076), .A1N(out[1]), .B0(n3042), .Y(n1397) );
  NAND2BXL U3370 ( .AN(n3046), .B(n3045), .Y(n3047) );
  OAI211XL U3371 ( .A0(n3050), .A1(n3049), .B0(n3048), .C0(n3047), .Y(n3073)
         );
  AOI22XL U3372 ( .A0(n3052), .A1(row_store[40]), .B0(n3051), .B1(
        row_store[16]), .Y(n3070) );
  AOI22XL U3373 ( .A0(n3054), .A1(row_store[12]), .B0(n3053), .B1(row_store[0]), .Y(n3069) );
  AOI22XL U3374 ( .A0(n3056), .A1(row_store[44]), .B0(n3055), .B1(
        row_store[32]), .Y(n3066) );
  AOI22XL U3375 ( .A0(n3058), .A1(row_store[4]), .B0(n3057), .B1(row_store[36]), .Y(n3065) );
  AOI22XL U3376 ( .A0(n3060), .A1(row_store[24]), .B0(n3059), .B1(
        row_store[28]), .Y(n3064) );
  AOI22XL U3377 ( .A0(n3062), .A1(row_store[8]), .B0(n3061), .B1(row_store[20]), .Y(n3063) );
  NAND4XL U3378 ( .A(n3070), .B(n3069), .C(n3068), .D(n3067), .Y(n3071) );
  OAI211XL U3379 ( .A0(n3074), .A1(n3073), .B0(n3072), .C0(n3071), .Y(n3075)
         );
  OAI2BB1XL U3380 ( .A0N(n3076), .A1N(out[0]), .B0(n3075), .Y(n1396) );
endmodule

