//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
iGfmSjTkktNQK5NQASuIatL0prK2CfujUsoKOgRMjpSXNNEmIP3SWMSEGN9XJ7Fy
GzaAlwSfZM++84ejceUfXDdy9PMTnwA3gsX5pPBbo4GLI+auIobf6QovE4kDsFUt
pQPjtDFRPlu9YGe9NI83mWjbud195/ohFwo1PyjZY2/pZGlw6uQ35A==
//pragma protect end_key_block
//pragma protect digest_block
N7f545O5AeouLByhpBGUZyli/fQ=
//pragma protect end_digest_block
//pragma protect data_block
/bNEYs80Vursd8URdxIsifDB5NOM/T13qjwrRDlm3EtdUp1DvirNTM6f2JPFgMe+
PVjvSaA5gdZtOWu48esea+s+AkY2+qEU0o4aKtdkaVJXCVYHe2uBQeIEpcibwJT3
V94/tTuf3H9Uu2QokwNDEGvTfE/G5Fm7eW21TKd/RcpwEZB13AU26eR4Ux2d0oii
m3RhzE5rF2spA8vLpQjOU3sq8SfjbOmg/Z3yAl4C0iY00c1aR4N8KEZZOOD7HwT+
xu2NGkyvQwqJXL2q2ACI3xs82snHkujVpPsAnrKaGxSf3gJ6//laBgCABESsHB9x
Fafy2yF5jye/V5GL5tLqWvzdd1kkAX1GnHui+2DPZ9nOkT5Fp9qUabmlu+SMa9dB
iNNZUSMcKY4i7dMBFVEjjRTuMCCPqAUkYbhF75MilUZL+5O9j5vGVpm+/OZ+7rXo
ObBK0NVWvyfWsyDsMdCll0OzVcWabQ1vwXq2h5UdEJcVo4IJ+00qmmWFuHoxCFTt
jg3//nQ7JdsdIMLJbeuC/hAEA+5J8FLoq9guCWuRKETXVwAAPpw3AA6Suy2IQcuc
BHXc1lVJFucv3wAkV0OovVZ86ax+GDurBNQIpe/xkGtdhYfuBbFFSyO+o2ltJzON
nw/4TIsV5H6LnEKTvwaCJPFlEp0NYOAJBfEQOihGCzQvrkrarYSsg9iA8uPLZLsk
rwq9I5rW0HwvrbOPWsGagi9L/LXKYkEAXZGvnB0/sGwTrw6CJPh+YVz5cFMSCr0R
fXuj5Dk3Kexfa3uz/VYlDFtRdkwA5/Djbj0CCJv0S5HR7hyozbnQtfbRpVgnlw6g
zkixxyeoPEuW/aFXAIDPBfCK2xb+RqqqeM27GQOxSwNDZZPXifAp4TOYiae2cSdC
TFKPLFmMawFFLgGjSdXuHc/GvtfhJVfK9WeRyuTdnQSd9wZMwsoGehkJ5DIuWdxQ
MDTeg16sa0FhIS2jFSHb7K00GYbv11Bw8jZaykldOQHwg0s6GfmZqks00UdO0xXQ
t4Sd+vJU11y4yBgf0WbWkj6Q7YTgcG2f6A+bs5PskMk4grRzOm0yg5INbND9SkZS
4lQ3/MxmbiAG99NlOW3Ular3qOapNpm36ur6LWQssfx4mlbQxuOdzDj1X54sawog
e0hnNRvhwKm1qYLk2G3NkPQVemynGy+/mOS5OveirodysH7FzzDw6EDPDxGGCYXq
ivL7U/a0iAnqZfnPaC0xO76WEySVJryh+zScNOgOkmgtKNJs8/N881IOrikLx1uZ
Luwvuzux7f84WZ/6Xc1+nHQt+QG2VhmhKW1QGVZy5A1RaR2OPDRRHzoPSXBIvdlq
/HIamwhQcRN37LOE6Zy20TBdLz5CuqNDm3QsXI48tikjxVLS146uGU3Kn1lyJKwc

//pragma protect end_data_block
//pragma protect digest_block
T+U0MTrjKqHf7UWEn80Mx+oo5MI=
//pragma protect end_digest_block
//pragma protect end_protected
`include "Usertype_PKG.sv"
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
F1iA9eW3STauXtvArakhsZqQf5MWf03JNKfDFuWVq2SUMN1bvtOncTiV2336lNAw
ykDirDeR22mcMDUWGcU9DoKNq4eBEVnH+ULC7n7vf3QgfCzcbzapHs3C3OOu02MT
bHuUdXSR/8EYvY4YGFWu+y89+cSQ+z+zaAZZ5ZsWzhYwSmBXULHKaA==
//pragma protect end_key_block
//pragma protect digest_block
ty0VEghrRoD3bm3EqpN228gtRmA=
//pragma protect end_digest_block
//pragma protect data_block
0i99e5aEGZkOfkNzSg/w4PRNRT8FXYhmoDVx7bOYMN2EMCViGlQEuWNoICzw7q3r
rhqWehaudYIXx6HH+qbB1L7uXg1+Jya1tnS5Ep1cyJPcyqXUlplnGPJthn2xiN+p
OgSxr0ynjhj2ol6ox4fHBM1pbWYtbP3P6MQ8svquaLB9YvmyY3yttW7EEEejcAFw
WidmEk349AF3YezXyusB0Ka663SYK8lnOTbcTMi6z6k0cE3lyZITXSvqqhsJzkrB
urbWEgyCisvPT46yqVe7Fds2WxzDmE2ReqzQV3FWSeOTZ5YSbJM4va3n59SUf+uF
h3tagLypMeqe8+ivXhiNgJpOTcgvNypDXML7u5WMbgqdQ7/Z96TJV2AQAyjyo6fH
JUEdvr6JOpxqeNyfCXuvX/jpNVpRfGtGOf6GKDyke2ySEXEs9fCD4rA+l0YzbM7P
kdpWOXy3YUc+C7BUx02nXP/UdXqnYt4CMc/AWBiLKXCsRlKCpfCNxMjuikvH0ttu
b9+mY/zSvgq/1CExz8R2PRXlRGg9N/hIcUaP3yz+oCceJ3eTI1hU7yLurqQCvSmR
bw2+76TaeH1Ki9emsKmym5XwKWYcLsA6LjuH7wgKA73INMBAfIT1DsvDZCyOkU1b
BCxgAYYrPf8vCGWXx5qT6+YcY/yduwYeYLVD+yum/ibo2ygtwRpT7z+YOJ/BbCa8
phH5gzSWotQxveZO3Ex4TEwfXMyQOi3eNgAqYFFjO9Dvweu2TAQBwgByqpEciC84
XHmyov6th7UP1k4gOQceWkiJpoK4Ng+ej8eIxgQ7SzghPnApffz/nI8E5bv4eOqf
i14uH6Aj2YAdNMya3YoP/rbkqIymp9OcWN8FfNfZMvqoiVfguDvrn5na/V1n2gdj
SJWRAOxdeXesyj+jvym2vfFZpKIOdaKIRHCGF+4Y3pLgZOjO3h5iedIUwd7XJWud
2gPSzcJJlbzIg2d34TLKxYNpSFrXm8PUMj+/X9Jp3HcRwHF2lnxFw1+3Ae2ZxFiA
bTCg/Xx31x3ZwC9/5PEyaIqg/1ZN5PVrhdYSzNEMm/Vt+Ub0qsmAraZgkwAT33Cv
Rd7HIeEA05LS76970qXlPmMZANxDQExlP/IJWXBU3EeGkuLSNjZQU/4rfkY5Q0VO
ACA4eW36+kgCkGpkf1UezR/8SlkTuQia5aPqJLfXHf+4pgwre5hJwdVApN1BU6Oq
JKwLdSgqrJZFNdfGpFAQS5IFz9xgaZ4HiH+fAieExC9MkxLYUHAmXTJTm3aJvMQo
9mxyaimNtZgFa/eWTw8bSlDwZHaVQAdLV58eUFL5W+k+/1IZvuEjNFhPx+ilWTrt
QrqscWfOH2KNt0T6fJaZ0o6RKVNiVjwf3mYFy0s8QZyXq2TXdtRwLdJ6TSkyuFEn
BjE2F4zUB8XJURN23OhU1jZVA4DvdwLqm++VvMsPOpkG2/WAOicjUIM9zuNr8fsS
uAxbrISOJOayGXlU7axfZh09npxugTzbJtZDiXv4CCh0X6SeSoZNhSrkiMpnc9U9
gE2OJOPNGYv14ghZBc3C9sxEsM7zRLpY51Nu/cszKqQS+8duv2aO5m0ARpHHz/NY
tFmU+f7Hzzl0bgqRBrwJ9ywz7KRXIqnnriiwiigxx87CaMsYlK1ZiC4KqHnRQ5aZ
hda6hK5I6A+ZfV2DrNw/Rx0gWdxGkzeVxIciF1j3/XpwdSDHYlLncq7BbsQrroD2
vX614pt2VhyBW0gh19jtwd4RPzUXXt9KSSDJsZwHRIA4mlKLEokTSkOkZytoAb9l
aBwC2oHU20iQHZCaGxoh/C2EQYFXmzCjm4eP8tUAFRTHYQjINCDOF5YpTnNWSxMK
6nAXvANJsiYnO1bThrIcIzhuK1KyQ73DH/hqkLxCmD/HKITi/NVWerQCcBdR62Jl
Jy4J2F6bzmYwq/SBj6smxOhdPjxQTibM6iRedf3GiIQwkrYyJwbi0wCjUBTKCr12
KV7BtrcCQY5trt7Jw9DIaLzJ6VmKfDZlZJm1hmkag7dov2PwraufPF3s68BIfc3S
SO6faazEyym7q45yfp2TGkI8SwfXYCDWQjLrBGhiwpJd2IV3PHYs1pTFb/mFHkro
+girLR6UaqyXDy7fHMh522P7pE+yd3V9S9/dJwIdtgyE/fcKaatTyb4Em2anhdrp
G0YaZXegsxN5j6ENn3kiJLF01lKpcad1oQHraafS4/If8JCVsYR1rMDhGVTRj5og
uLZzbWjST96CNTCCguFq4+g3TJ7AAvtc30kogrzKVgtRtYlGlss3sCpDkzLrgC0X
nqME8cJwIVbLeK+uDpkDBZIEXpCwGO/CghZFQHdU+u3e0oBexvveB2lWoi5gWSDz
b38A2r8/t5iPFajAgacUq3DALnOc9z4+H50lvfNe7IZn8l7l3+jSYnevM5Ro9RQZ
hotK5t/lzW173g8p6kZahPWnWaUAbZR6XrZq3RJanOzoe9dOWxzKVIlGnH3gWDaP
3Cyu5BvpjjGrqsrdSxzIwW+gKRiWodCINSF0INx0yrm7XnB3X4o3OPNLXvVotHLx
6PwnP+kW7AZe+KYnOV4Ki/vTa/niu35S+quPeHoFzLA0YneYS/7kqIshJ/mMFEnc
XE/3RlYv5x/FwP31lFnPDPjagGqyT7/yO0haya/Qd+y+8akPOrBYSHAQKLtHveUM
kVIcS6gph6dJytIXt1gnDdF0+IuTirg3Eo+Ch09tmV9vPnMhj9RWE9lwPiFkHYE+
JLklHTWuvyLKleWYj6MZ21Cpqhm1oNd+hwRcJOb8cwTSYbuhkky3bA1OGeBzQXxi
tr4jpFjGTKume7BNfkmkDA0ET+t7tR+siP9yojItL/ObQbVI4pKSaBtesU1wuBmQ
N2e4CwqXtsdHYrjqy7VxyyLKHL9YwvzfptlHu9GJtLttFPcm8FKFIGd7EgcWt8EU
MrwfuB6ezYibUWcEyaXtKLm2DOEofT4zz2iNI+JNJERVzTFTVhrmdWJEPMTzILz7
su6dbbZp9z1Ix3Zhy0r7LFerAQ6P/aWXYK5MCMQQTgVvW+FLTIqGJC6iIYE85psA
J9MhHRlioBz/UipCk2XTxrV1LnyrG7OcpLpC9UU+yI7VG2z4bMy9V/uWLVg5H/vC
x8IeAYO/1O//1+GphvwvAQFXZn/G0Tr2GpnVHlD/OaJHL4J2UzFBUm3uYcdoYy2h
tV4nRy+TqYhrgfpt9FMDcQjMyptINPHo9uURxHg5MhAoyn9utlwvyzmIPlqjkDyT
Jqx7dh+6DgbdLiKRA3Gnt0vwTq3VJ6I34QoDlutc9lSk6GJhqJ5Bib8oeS0vbYo5
t4ghE0d8tPxKI2MPf96+ZENeXtakl76iPasq6mDUggiByqt6Vdd+T+kvnfihyRSH
/1AeHYc9vDf/e8EBLgW97DQz3IeQN7lVVZ2EkBC7ZgnQ4Cah3wx2LNCRWUAQBXUj
+vl1eCNGI+rNo+Pl+p1e2jyeg7WByRmL9HRksN0caRwYrI3SYO1eCinlda4C3Eq0
P5or9aKRHPpIUf+H55h+OZ7TfSMkyxv1mRVGkqVpjJXT+2Shohe6aF8tcTGa1bCx
4tOQNrcri6YOLCU3RX30Hx1fnKD1t6vNwtfTEGNa5cWUvO4ryxkpzP4FGznuieKW
JpYvMTdm85zr5FlNQS9IUub6Rdp3Lk8vV5/C/ZXoACZuPI81yycaicpDTggIlVHh
Dqqjl7GtZKefQCWVpT7YWw435ylx1zt0godtz6KmFPaAKheBCPBYWF+JZeOPpVyN
JUys4OurreWh9YF2mgPbAbIMrqYcpr8U9H5aYfpdzEaQPexVXSw1n/lrvTj8dBTI
8u2RzTpXRhnwM6R9M+uqvPucPaLG7LMbAIIBgx6F9/DFfV29OmhwDjZQ/szU1UTR
KrgUc22T+Nd+do6SKd1EONImlfjDd1vy5mih7s4HwSPsYbcir0YF9UMhaDrjLY8D
HpUb8lLCDvdEazs/7zmT5RDO3IB2Rrj6jcR46D00tsJfG4AD5ntjRPfe07hZgenA
G3lKn0D2tu7xzkioha5xS5Nuk6ife75/abtdeJzT8n4VeGbpgt/3Q/6EiV9DB4mm
4Rs94NfnswUpCPTB4ST6DiCNaHXjsaUp9E9BOKpBLokXqCRwmBfMcJSFTdovTZb+
Gzsu1Qt2kd7Gv6Ubf4oqYcOkkfi89Y0AATqlxzuf7MbNL5FvK5e23u+bVbI2SXbu
Bst6T7gLeAmGTavTymJixO8PcKNLWLcRAqbrmay2z7cp63OG7rypt8kcsH7C+0pt
2/cCIUMjP5bdDpjLinwsq/SWwPO198VOZj+0ST4gF5UGCUfvcCG6rY8bwxw2FvmX
hWp2h1OjhL4Muz9KzWML+Q+fGYjuClnzpzwrEwBIpH3uYuollUpen7q++YMHE+JZ
4f94O7l9tpieLkqeXZLlfFtnKAAt6XXAOrnj5WbHU9PrPAzQs+RJLfgiFzG7OoGT
Bo2QXZ0oktY5nTwi4oTFPZSNkUoL8Wn7J+rCH/LgHSerz0d+dOG16mxzBLPLlAbP
DWiNcd+YMFJCSj52nqGHzkGQWQGS6hKIlUk5LgmGKUZinWij5mKv9aI3b7r8Jkl/
u4mzwT/JAzgsHjWaY2CWZJMd8Cw6XeYnYZbAxS6BgdACCv8PKu60baHSd57+JLVd
AfM6AwmaztXt6Kxk3UQNT4Ss0O883jXKbnp1fiNTyaHHSNtNT6qUGUUUZRGznHpZ
KfIeXSe2YEVyJKMvLFecnc/Pm9wpka7jUtg0cYqEcJvKDB8+yeEDaXqlmelja2bR
5/UleD0rm2YZl8saMYeySBTx/p+H/d6qrVY3W+EoRpLYgZD9YOtHAVySaItPa4Ih
PvHbMqF2FQ3/jxWlxBM9DpultxJHNKbHYfo9ua1TBylG7WyScUlJ3tJ51C3VJc8x
nqCZL53KzwrWcC8g73QuR+vkVHnAaMXwSweNyMQs4uyeIhuBRWEH3AFcLGF1aLQK
CcGz9zNP1eIm+J5B63q28wwzKovyX0X50y50M7k5eDg1xAXYl2oJjdDpCAnh8oB0
j5PPs1hT/jtjPFnd1+PXRklKsffQrtolXz3sIP9ZycKAHzqcGyVL9Uvt7c/WU+Gn
/+JR6uicx3Y4dDKMFeyhdsPlEjELykQEMevKk29wCF4ifJe9AoyNgnyQR6KvIm8t
yEXmcIVO63WITeFa3kpBeCBLQQS9nG1bDjuFuKZbS4hthSKPxeWN1ZK6Rghu7e+z
TRyk+1tc8PrtSg0tZ0CE81nH1hpQuFA/o/dgYlazssCjjoPqtELjRLph88NiHj4X
276qKSHMugQ/9xVipVZdUifjjKhnPV5aPUyM+LYoeL37/w3AfwVQB7IQvzOS1lGm
OKQgZDWAPotpNVUWdexb9IIaJAUE8Nj5NaYUlMTni8IMtfietKFR6DuN/55vuxb4
b6tGINJRPJZxbHFlIx34X1+fSNteqcleDawu4V02DEhPfTp7LVcQ/IpzbrEvYlnr
aFS9dVAlfb6qwdpis5iyBEpdhqrBONR6niqFCNWEh0aYdY4Uaucpb1exVcoEIsRb
Rx8nKKSpptndV4PUVdLWL+CaJ4ci15zDjgVXsr5QzkEenZmbFOkx6BtqAxlxKQ52
2BBSxz4BrFfk9nWBau/ykt5ZkoPIQVhTRlStmflewwQlZICBj94bRz/fIt2nwk0r
Pd3/fj92tWTHJJ4HbS/YBsSJzuyLIkC/waXvSKUos0iJbXxi2bS2j6X9NIcAN9Wx
gHX9hgHCRNS7skVOnr5O8SyWfLVILB+x1wCWp4eCb4viWQx2ByUy/klqMgEpnNix
0tFhbtGpGmWR+xTqtrpLQkril3LZ6hgI2WXfjOgVUA1fw2rorqyWkxcRaLM1jzaP
uJreqy+lDSA7nMD3ORERfYM7H5dcVx7ol6C5qcWG5IXF76PyLfXzi7trUazSZzeD
AUBL+A8ffISFob+gLqmrZpZlELjZ/cyqePFwzkgTSqGbVxc8Sg59k3jZ0YLHwS0x
nyTg1gVqM0pHVGTUzSOVHD+P6qq66kfFptFD4t2eRoL9JpKgkg3us4hF9SgWrG1x
9/5DCKv/2Q+PWAYuAjLIJZS/V0e5Bm3X/YVi3rHRVnakVLYgaPYhm8vq4O6gECPI
HSehr8YPNHjK/6AXYublDpzAZD8+xSe6mb+SQORJ+ps1+PiGhWf88C7JgwnkPCCb
/uKFYCp9iRCmYoU4hzbQ1DSzYGFspe/agF/yTl4duYo+AkrQykZja+rE52k7Niyn
Kv/5EGqYb0vW4lB6MkbV8ax4QBTPujNj64LHyQZh9JuW0f86sKDkRvce98s3WiMK
3MdAaDhJMYEYg9fxtdMozXCC2XKp6V+wL7miKPv5Ahcrc6xSmStdsC0cApgrobvu
Lnml/1VNqoPi7KlK83xGpW/8Qj/gc4gC6xtvm9Bq6lLX/haWI0mrK/epQYJU9seJ
4q7Gl2/uuw/ZYlEEBU4mXhzQVHPRBBuB/6reprrIJ0iSyuNuBQFiRpTEe2l+9W70
wS+lni00igRmGRD8t1l7a0vEZ31OOpPK/PSqVo9ZadCZzrQkMdTFFhQSxrZ0coeY
gtFPObOZI+W5ACbiMsr0E5e/jHm7HRjAE2EpqMUndh6kxgw7P79jkn68XiE8a1QE
ttT+n5+FMGYTZZ5DRNekTQHHaVhavpjP0y5ZMNIGtsp3EPp5C31yxRYfNEYfX3P2
OuychpphBajFkJC+PSgBVrGho/u63F064oS1aIEPepZW+xFhQkI0Ey4dCPE03G7P
wT+GYOWKMQNnk6PfOe7GYPV8dcoxNsZi9/p1uKRSKakPiBjh59B/VcIQSKggFKL7
Y9xQwPaEwUvJlrXucYWVRTi8G4CZk9ypQkcrTqlqMDd/hz6sRQINIAyqDYmpfVq/
5a1vGSgTe4QM3qwpRIApPXzOPlkH6mf/Htyt5edDd6B12X9JZbZjK1aVIP9nUqUO
kf4/R67cCSBqCK0Brq1h6Rxvp9GRytHMtSSMCKLCeRhNK8PpDSxT2KdEzyR6X6f3
8ln3OGFHe6/DTagSUniIQtHdnbVQLzb5Xi2Lxv8Ad8v5yWKazr2H/TlP0PTLGQ7L
X+OUSqe9z9PKWLvvJQWk5EqX0X227eUJED414tEIOzfUyRMy0tTIt7O4vC4cid6v
xKi9hFfvmFp7lWeXTEhoW1q+/MhbXOZqoaYQPVlhDLxJk6fg7zCEF2W3Ofxsgu4U
cUG7BVfw9HAI7OfmNl88ZJDlZB5x8ROqNeE6BjbGpzA/rVCj3Mx4aKnKprHSS7+Z
kDk2zCPhQwzRQA8OI1cr6cAkLIIHAr6pcCw+u2BgpdcUmsCPnl1ewcVEuGNQQCH6
ljPjKdMY8+FpMc9qUjZetzqGms5SQwyj7RcZNS1sHCj3gFyYl8X0z1n9bFU79k5K
OJotL2IaDizvN/22ur+9E1lLyTZg5SuCTZYlxJigQ82Uafd5VqH0AvBogPtXmqGy
QMu4Duh3avg/e741zUt6j+Vjwh8fNBgHTRUTrBSIFX6f0zhm2deULwOihrxjYsZC
Zmiv6kB6djBM1kx/DDEt3ivDcFIw95OyItjcYHhx1+CYAIIfICYVVA97+6bn9Hl5
VjSSYyQF3Rxi2cQHtzhgH/fk2sQaYx36AS/DX1cT4MLzXfkS2kgrWUjVDjAvL5aY
8rIMXUdIe9Jn2fqQdr5VjzeIz05TtId4D96zEwMsimb0qRd4+RnSxwEEJKcvX9qI
NdMEezGpmsPqgEJD1zwiy1+Or1V0zIaAKn9yS9FsJeXNNC2XIlTJEd5UgvTCQn58
vhBbdS7NNbIEGsHZhx8Ljzn54jqDNIXg62Mo8BE0KtPGI7JsGGfol8g9+4U+V24h
IqUFMsft2Xv1T+WbfpXiYhHMI3UioouPEROiMHfFDUQnUQpzFP8YaTxBk5NFmo0J
1agQjL5UPQJdjlBlBeP1aTF2vWdlHe73JUtd6oqyt/N99m7em0JdehzRAVrH5ljI
KFhUEVQB/J6MjJh7Ma4uQDvEh8i2xqYMQR6eDPms+2m2Y1cIsWMoCnYxLJRzJnpx
62hIHHQNInEaRRztRjOkZ//m7c9ixMe28uvFJ2wEhCTyGBKS+6NSvB3AIhd6rE4L
yXY1bG/EOuKp0R3c6B8fD98o0XK7mPRLK6YCRKEPGOPdz+ELHzs4DICt9CkCvrLi
DgLQjgA3sGUenwDIsgq7EKehF+2K1mfxkSqF/o+ZN7EVSHPY2ZEVc6PRLeW+tZux
1xmO1rAyRjwvD6dfQV95VKdSM+qKyI6Irxri/dhNJJ+xSOp498GrCr+FqP6y9xnt
Ii3zjiJEaFzCBoPfrvP3pGm8yEF33bDwGc0LsUVK7z8KPPg2eBMZfFkukNMU1uDq
5xVyQqUcECIcljgXdx/LooRoookO0eq+QpJVvTBuYr4R4ZTCmFovEXK5Fx+s3ZBF
JWpb3tqQ+uizgQaow1Wn13QjD3d0ADjKIIz0gpgONbjaZQr86C3sPhM3O04YlEs/
hjZNKMKdtECqRaxQvxYFnA7iWAat8332Ts2AffG6XTKvKesDl/3KixOKJyAfbTkT
HYZpZhnYdwu63Fjp4CGnfk2AjbE2oWi/XDZP8yL/iq62YCUyiARwEbcUOI3kuDcW
krxBJSmDmYkTYGKMfTcB4Zn2MeuRo6LKJ7zbvtfqADvna5iQmhDM1wcOlO3qSZMR
RtToPT1+Vbyp/yP7uH3P6/zjZ/jL6Ej8cVVL0Yp1yufTXBCx4Kmdq10uDKjbTxa3
mb9aXrWuh2lcxRJy37bS19QCVymYFhr99e+8U1UVxPklwceleWAoMYAF1HX98Uqh
N22Q7R0sNDVl0s73fm8QCyzIIMBp9k2PB7EshVu5V2oRDu9B004oTGhl+QyYcRQi
fvbfQZ4G0Z8k91GV2dQuiMDXlHxYTwkPMJNgYQD5rR7o2T/g1QmFYCahWCPkxJHb
r+pWbL8I/XOG4MutxOd+fSeuTElBgqWY8gjAoC9l4QeJr11iODB6kZr3vIzPoAhN
jVoWfEeLQTnHM0iN5oXQQPdJlpgN5omvuhCqnkBH8GL9NQWdzDGpl7UpUJRpBL2J
aOkkczEAr2sd6QDT9Kjvrx/Gm9dpMh+vl3RtjSOosXqUhuT1XuUU7X2aNfZe+vft
v+mLdDb8Ty7jjLcUnT0aX77+YC7F22nmPy+n3MG5qv0Zb0wGuS85UdBuQBK+CgL4
AZohWycJYTwTnyG8bCoOhXtTMG9r8i5mAzIY5ahoW+lnIgu6vBI6FYZmiVl5OC1h
hcfVWGASXblYvYpA+8tpTTBmUAU3bMKMLUL0dhcnlq+WdD4NC6hPwhosZdRlVmVk
7v6FDGLQai3GGyCrbdU74WO5NJtebg/os6wIDm3pyr8ygkG+rNYPszBRFdwIPdI2
diKtVrq8IfpFntvh5rxuVdnA7IWaSmhFxi0qW6b+6uCT5uq4CP3E8Tukmxuv+snd
zMues5GKH6+HSNO7M5UVpy4gJX02HZwIuZXNtLIoqBFSiHub0JpnxmBC97zqPcdi
JNFyAoO7Otak+ky2HbH/LOcEmhHetSJyBEIhCr+0oAMJBYj/R4z4L4LAlP95XBn5
Qg4PVUJo4JyJlV0liX8Sniid8gGacZ3iErZ1LWgaAo0ElA6WV0HG7IP2bn8PMvos
KAei2WGg524aqbcivSGOVSGD1wBzRFGPl1d2FfpGinJuhC++RA7035A9MUPpB6yT
yx4ZENI9VxiutBLSNo8yPMeYnnSc5NegeDrnVYcG8X/Pk14tPUatN19lZCMWgsxV
k8a6W6SXWI3/RYCGcwbFs+JWf+n27bgwH7pJo1sdwtgG/y9K63q182gFtCdxL1lM
G7B6+o7V5Duj0aaXlsF8+ToNpt4QMEjTCIU/X6koOA+iY5AicEEOvuOjp5v0aiOH
Mml59omw81ca5Bm3tcIUhRnNaQcQ71+VHV5OPvyV/UlFDz04SNJHyOYu6ghfPOkV
a/qVDtIgYofRK5whWIDvkHMIrSD8H048G4iq0jMrxuRLB4Tudg8y40TVXgwgN2L5
0u2FBG3bL/7oUDrof2O0wFML5ueWSIOlakbYWJ4cKZuYu7r7kLhh8ik/0F3ulkyE
wFJVV54uNyZtiaioq98wRMd+ZgC8Ua3wFc9qBgzaY2+/HTAKyE90KdzODAsyX7sr
t+zT/EsVN8B2RINrNYYONpltZUhYlWdLg7vQdCZbxAvP613YAUM5dSqaf288HO40
uhzYZCotaShgblVj7qBZ/1i2qT9kDrnJNUPWw3FgXKx8gN55VKYpeG4Cny4Ul1/K
RbIBdBDPrI1RYv2vLx9UlEcxY40xMq1DaM56BNB5CYrasRhW7tnglLFP33Ek9XFi
+Bmb3tWFOhFs9pd6EzTn5SbZCdc2e3TSMrfZwm0Dq7RNNkzDFxdu8SxNj74OMMIL
kODZNOsEUeQEreWbUMM8vgx0pGLEvYKtnVXinKxpDf33BMYtOVkxsJRnyH9wOHgi
2rsatt7k0uPpSwhOCkWpbHIGOHOEfuwyC2H/IGCYNq6tFnO+6Iz//FsbCT6Fqo0t
+jmjyplRqutbAjcdWXQObJJOJynwhrlZ8UyTgDGrcWZxtNW4oY6tt236qH7uBdtU
7eVBkHLL6NR5rW9CN7hdvvwgA9azg700YqUSgW7vsVIOF02KpCyu0A9n0f6frU+E
uUEbZjCksOCuHxWJeBiCo1J2pQZB82H1fNQ0lEmseDfIC0UNYv9oFS0ExWkweEYk
pHOtkrdzVywxxh6f6FITwNySLmJs7dW8uDnQQAA2/0iJ0C1sW+6ucmDQaagFOvFS
Nt6TC9GGiINYucjDALsOJ0hpkqcMAyruneLjPQStlBt1K39ZanCzXxe5Wwd28t/N
IdPCta7ScjIVqbTUb3pcak93ejTsWATI+AJGbYUWW0B6ZWxwpBPhP2mng+LLzHzv
Wvzi66qX/cZcUkihrv7/66H8gtFfiPpgiCP0230Bp6LAvxWcKkFuT/KGcmzNDSOY
G2IBsMnFCwx6BN6O0Y8ZFfAI/sz7eXQk4GQ88L6uPKaHNApprua/oX6C2ULbLgxU
2pUMiqwR/tC7gJJ9U/mYq57T7GXK6qwDMx6nafSBoRvljFgv6afGz+JXZUD/r2bB
TufaYIsAEGkb0PGKWSJ24nB3LW/PJRfKc6tJG6G5tR12X9D1U04Vm3FC5WD1HGux
FQXkLkeSSdEFlz8Kq5XjUFKKJD+qRZe1nycF9XmYTU1R47fzFrs7w6CNznUbueO9
7X4k1FT7ji60tQ1hMPfnRsfCy2JsaoN+jCs/dHve3n1LWdmrDsPwxiw3S8yo/5nJ
fiQW4UcGNedQsWbdAphkJT3dho7ideYgVaNybVPG1yZUfDPe48I709b+NTPLUC6e
mbqE6UYV2lx7uUeIs3YAjNbUM2FKDZufbgSQ5g9FEmTUg+ZPsmsr5cLmyk2yGPuU
fwjOSM1g8P8uZoGknW1LxqXj+iIvXEzKPmsJCF+vRT73Q9TIABDtnVB+CJvUmz56
XslFlZaxDbVlB7M+krbB6jq6DELq/xnB5qATw6Zlsq0eVhvhldzn9ltB2vVRSQLR
nKuDWPF5qIbsl0aAhdxZahc3tOnd/9FjyPN0pd7LPIBQp68AGXMAbIbX/i6pjsJk
571yZjHSZeL3qZiO8p0ldILJ7uzXPabcUydYW1edgBn/OyHnV81uX0yUFh+x8Q3J
J7avRcOYV0dgyPza/E2q3se/EKyBDPOZy1zvadl4mWbTkEFf8hOyxADioekGXLEC
lPLXPC/iiE3mO4QUzMJ95orER1BXUzJAZXDg4SqFlyZC5nZwRqNZXEFBgwyl0tyu
QF6zPC8jMdvmoAyFNVk8PF30Jg3ql4IYdyA74HqDGiV/UmRKsMnmEd8Dp+Bno9Us
Oljy3jHxOgNibv1haCqOsWycdwfMz4LNXPowNFPZ8958n49axElVwQ2ivy6LkOvx
YnIL4xWDN+RiwMaMpIGO+Oe5p+ICzpZO1ZsGUd3L9NG7IdZHRVvhnlB0hI5F6x0y
Q5yQqkV7xqWe6M0Xpg9s9IvT5FwDrCDGV/brKuoOY2r+ZUkmAzJeiPosMdIeHD8m
SDblq8zeYrnc5ER15KF599qeW4nc3TdWoteGQwy3/M3f8AtY1/jE1BfHyy6Mv5T2
3+CT/S+MJuMd1aT2S7Op4dPNGaol08/LpclAV/bGWLVHo2KMOX2iZSJZXDKrcBgg
JiMoKGCXZW+XzjBYCZt9VnvAL1lbN9IHBDs6tzOZp9Mgb+UAgtwNE1PZ+5lwJSPz
+eJXRP7vzfZkcWbp8QraYaK9JqKHwng8gLRyJLFmJ98EQ9+tYjq+X+O10fPFbv2z
oJYCb3fmhSy8xsK7aE4F88k1S+i9m6aX317zVj2MBVyuzpbNClyIWsJR8DEBWVpc
xsxS9S7USfpK+CiWXAEti/gE/DVNycnu1bxT6YjHrSTdaI/0B1ULWUraJdk/cT+S
wB2ow0nDzisWgAkGF1XvkLXIwiKw6ekSDrkJp40XMyPTqEh8eEIT/P8D/BRFd+xF
iheKIgOjEYruXgJR085d8osAdmfwuB0/608RktWhaA5Mb56K0TuTLy1gZ+lT1GBO
ECDipPHSIzj70a9FDFfcvcvkgAdpU99NHCodW8TLWa7EBYGNtIKZrpglYd1WyHfu
4+dJZRWgxSOH9khmF926FlYetCr1m7O2MGMRutn2dFUFy9Lw3axn1KSAZmmpQlXd
r8wriORqvm/kPrPn7XNJAIGcMNKk8WKkjzGP5kvdmDfSocjTnWp0xJsv01hRMMqp
XVfV3QXhmziRUNxiPgLWLOI3ixjlCI2GHMSW/4E7wtcZeTj9z80b/8HngLscHwZ8
RV9/A7LT0Jx0EafCy7MBN4BicuHnR1OgtqW2hTPGSaMIydogB7z3LvF45TcrWYBY
6mW0Yr7mEnBFymPX4YMhtEdTdhzASTn+9wjOTyRTsHBbfhvszWPBwiLQAsSooVUR
u+tU6QsudINfPFDc9hnmkmhPW3nX3mTb01l6YYB+GiK7ZFLmdus1ZQCoH/2hbue0
Q6KCY/WNNFxUxNLvhe5oHJqHHeFEB8nsbynD503kgbgLoMIUEmBUzNsEnkDA/447
/los4Oh2o033ZZYdVvceU+5Ht7jMTVJzcoM9kdOtz3uf4y2T5E7Ar+ZtVsDS2TiM
72Od+UNKTjzjVwo6AuF3TSRa+FWEOueuuiTCJ7s5TpEpX+E9ajghwxSg9rysUFg/
MP61CxD79hwZqVhGU0Sm/32N0EtOiKU5RLzWE348QRG3tV1EwW6mrx6s2lhEc9Fn
mVcCISXCIdeKwazFyenhR53cEHFAjHhSDgAEItc9VRdR4zg5aNkPoQHxII/NerHq
VDSLaQZR5Tjxy/1Kbf8vGtNcI1dSwjpastTzIijVUugq+vqeo2U09azmmJd6q7FP
GO5nXuKiWGZzJhriyOxfXUaJ0FyFoXLwRdzHmLjirpO2cFHa3IDp3ZK1+J0ljEvp
EzPschoEZOgfWU2JTAZMbsMxvPBTh6IrCRJ5KA/ahgw72XLr3hH/UuNRx/+J8W1b
4KFgqA78GbNkyyWsmo6IV/hGK1HUWPqEHHfJCJuFIPil0GwfwopLSM18bHNSHK/w
AAnsQWAZJyNHiwA9XtG6b34NiqPabnEPAudu8pdmh1BKu5NU15w5aRrNyptAx9bW
99Celji2+0o8ix7k2e3rbJo4aMHurXZADwTpzJ4j9yJIuMFWGH0mgVkCyJnLd7LC
JZKANykVy7rnLdSpE9lMqHsrMsn2ZlzpMMYfY/N3yNRRexFYf8Kq1TYwWyLttRg9
Tsps3UyktxXSJSX8Rm/ennNBCoxicPbd219i0B50PEaJeqjelVZXRJ1mKR7SRRzb
oJSvbIhQobCZj2Tlj96OWCV2QZBoSykRjsGen/ODDHKhUOXqms2gXRDxIvRJJ2u3
XVdlEMk6O/GevO0KSu4OfY18xGahAozXf+XCCO6WKxzdFtk6Th1YIvcRzY1HZupm
nFxW/iX9MyEChL4hWBrHwOg/1P61DBq427L4W6mEC/vALcubLGc3Q6TQlbQCyVEv
aGeDC/GNjP+sZlH+xxIXUb4xDd0AJDoNlB92A5Cu7Ih/Dv79hgwRZWEn5OBrWPd8
HIk51A5ldb3o2Pd75YL3zBEg9yJorXohCx6bzMqGybmJYtvJ5logrYcjtkj9Ey35
h6cfkjV7OK+9l/oSAtZzly44EWLKrqFcdw3KGgnKv8BKbVG09AbbknupY+Hp1PeL
Y8zWenZzLV0ZVHUERVrhjHq0U3pfHz8rtRl59dWkydI8hPm8zBxTLPPx26Rj6IMq
e9QhevxLy0RkQmd1DL0mTxlsFSgIli3oC5hj9OBMcC8HBTbY/NQHJOzrrS2IxsBC
SquOAX8EfyKIEoAt4e7yum0w0c57D+13qbcJTk/RU+MLIQ+kOFR6Ixo+oqG05aum
UYr9xRadQ8eBVoYiCbbifI+4a+4OdaX3uf/qiHKz6dYXNv9yIOuNknRVpGKPT6Ol
yYcTNc24nncmrxiINtZOalqWdoOCupfPnX8b/KMEgfz7vVA2e/ZUvKDJrhtzwz3L
9GwRc4nNvbBRDiMcyDuvcRJK0ptT8hrL/ekWzu0IaBKomqNSL8vCfUrx42y+e1fA
1HVj6hjbfxJt2j93iL9cSV/2yAqlIPYRKjtzjmalwJzgjX82TQmgUaVac+CRiSGq
R8FmkspJXDB5qivrrkpg+mwA0J3gzfcvb7xM6HD1oTzFP2HFfLCd9JYFA4ELtxZl
XPYnNUqeLnJIu7AeDz0S2pZZnBEYqTRO33bFLrQRRDVGlmgm0g818ArimuFw6Tl+
OMkKL5QfPpk1GaODV1c64QkQRGoHpBa917Soi7p+QBJwqGmJCxWoarS8/KtSt9pW
fwZ+brfbNY7jbsb5FhhJy162Rx5Q1j0B/wjXSC3t33UHaRxRdVYBtcUHN4XzpZz8
pp2mfT+ciS8MHd1gHl3WoV+T9RwLq5dL2RfojVdVjPkglhKZiMjN2l41UYJ1bhG6
VHPHUJQatJLMnzO4KzOl77fqm2kXX/GsIfRCwHBzSn2xbL6jsRsK1cu8B0IS7/dm
Q2NTITY9xjKVy0HnLV10HMUkO/mcHjfxaqGJw5JbAJuEgH4ED2HQB5+2qvcpDXFV
te6PF+bF9njTjdF51ApDA6VaGaiv4pWUuEdnxHXeHvW6wKIlo78BzWYDT9YuJ7ZG
DYD3vKooMl/LR0zvsFyNM0S3tQ4HcPzTABTUq9Szr8FPCpKJOn6wSOV9lehDf/7a
vA1/NWG5C1riqJXdId7xRYu8BpjVVo1w3Whjmv1SYNI+oSVMNWeClfr0+U+nz70G
8DmyXzZ4/Kp/z+UbOBmvVxFGfjDd4GLmrJstM8UI6wLSOevmWUffNFZuqrgimRfQ
kwSeN7lfqs8ba/zgpJ+aMcGs7Js/qj1Ce3KbxlUr+cpuzTi6NPH2ctSe6nxEXOS9
qoJdX9mhuaPX3+hkj0YIsPwBWhvIidhWRvLpI6Lag/KVHRWsniNApjQe8k3YX65k
S+i+cv6eFlXbBJS5/XX25IEB4tn3+/QHXgBYYOczu/W2LRjDV9RXciRQfJJnVJ+h
3rT291GPFsbjuB1FGlXCrUk/uSXlyn10u7Zi658Exma2D6bMYOG9I0di9QP6NiSs
EzYCaSi3lLKoqjS+xZGqbZowRW+3u+uXeJ5IhAKwcAzyKEkowz8opOnhTMNmPRHp
KHwO5s/F3hEXoimzfyGCpD+CTERxSZBHpzSkXFMXaAcCDr5uMWJtkqnVKnVsgnrR
e7stPxm5n3Vq5b/0xoaLXJlDzGVBRMpi4DsXxcMdXy21dKqyJSB/zsNnVWROeo48
I65HikzP/4BQ1cpQnb0UwjiHdtJrbXpeAXxa4KE1ZiHVB5B2G6DjTER30s9rJrxA
UUZhJZfF+76rvtfXhiqno27dlfOkmUGpMsflRPZhGLqeVQIXBK7vjr3lvEgCmAS7
DneABb83BzQtd2in8BU9PYfWGhOwosVriID9pREibiwu9FJ4cj/b/AHqsn9jf9Ai
bCbyoWaq9Z4ohSM1sH063jUjg7GHaU+/Emm8XFX8MfJRkcfehGYKXnUV0QP51A+H
G3PdO+VcEsIpJalTR+AXzrLZcrzVA3Rhgc7E0A1VnyYPkqVmYiC1dO1aknY4LBjF
fZSDBaium+rhBDKvXYXzHh+D9ZXoBtkSgUiCLyR5tREAwrdHFw/UPk41UfbIIRKh
XgpwNjMQ+gmmHOITnBySpfNo5VUreRymnNpXD/ot/R5CLtYmpFwfiaest9ejpk5P
mrzs6QRcMu4KBct7/2jCa2lUCdIkBKUzJzMgfRvw5Zpbtz7bQuCGbpsKbudNYz92
J5XqDqvSJdIwv+Sa2Gs2uchESngekpuHmyKlMlSwNEX4CSEdn0yy2UDZEYhgyk6L
5WedN1aWhjDDiwhC5py3aSvV9+FH8OIEBMaNl3gAFqqOY2ESnbS3X60dwUMFNGKA
6se7+LJJAdJQ2p8UJdruiHMrU0tWg7aG0mcSxp2pLue8y61lZmtgG1zd8O54Vmzy
jH5u5xsIBsf1jra6nDjxgrjiDyeHeoFKB2dbkIRSWeOrPESzevWd26aSGGEQxXs6
mIfKxF5dBWsBMAeCw6JFi1l7smiHdE+qNM86keDYAKF6Clgaf43uXHpifW6kARO/
knB542rZlW0RDA3UUmxBaHFNH3pHhVOBtgZjgK8JCjUvBLh+pGA8hyxTV1TFwQxb
y5+FqUGvCxYTI7My2sDKEF8Fn18oMYJdtVn4dDq6gJptaCjeX5cGmVS/LJWI1OsY
f+6jNzjhQwpIQsoJJ2f13i9RfginRB49X2eCHHHYfZFbYcJNmqgdW9to9/vsHz7p
pZBk274FhiKfpsxpjtBmBucttGjvPnbfNErBNcXFFoBrrqaCgKT1inn4rVP7JQLA
N8JMThe/1v5qNl/6SVmfCU2tfrdkuwy9hbM5V21BQ+fLsgItxj++d5YRxqUAndP3
UclRXz2N5ko4Oivt4drwbV+u5wnJsj3GKcjAdOrB0HI1iIFgKYlxHP9Lm4sUtWBm
jSMpziTFFEPyGMrPbFgqvu3dfsviC86HL90WK8XK7d9qUHJbsIvk9bqhRLwUXh0z
gd74N7dU3ZoyPXZKrVyaMpNKC2kCa3x8lK5OEYQq+YJcqfSvk4HjGL3dtO5mdQtI
gcnYt6+Sos1OPnFBqZsE1/ouf5IVspX1sy8A+0XD69WrCHZ7sY+4eZ8mmvqcoU4e
RZ5nnbFmHFOW5ve/U2EWvb/y0svFAOe6G7A02OnZKgfNS9G3Ieq1j2Wa4XfHU4tJ
jqi169r63ap6mv+eTlORtGNzhdENJOS2imOPF81j7RV53GHvb4rjdIM66r5t1jJM
eD3ZWgoziDFJC1Gpovw7WCC+3bqJ4p8TMpNEypviqZ3sMUNoyIdgCQFMFD2Ay7s+
M9fqYuMkSdxXiPTRAEMTADMCnrOYPCnCWhoZBDX6fWbLHpkZ7OUJc5hc2GsOqRrX
DjQyW7yZP0e254DCdLF+BGXt1zIFnl+FI/RkJ6S/QYVlY9dTDNlaCNqApjoFu1On
8/o/CyuIu5rMI0bZ+DX17VzdB1STsLK7Q5crLXIM1CHUzqhYttFVb3Aucs6yjK3o
VmPkGuoBEAk7K/yRzpCBph7Ign2ExsXG7JR6k+eG+i586n0FjXgu6obxufF4FXSb
4+LDfwG7ZcQm0J4tBhmuzahWI2Y6Sar3GUhMoHeTnp3ihV3HKkDGNgnkEow2/mqR
ToMcRKDtteailrk+UMv2un+mGHEJ7WgSi/AeEG6QHHYiIkwo3O9G3DCg+D560TOF
/qa4QbBjphVyrta59cdjumpR/6IaJvj+QfU0ua9GtRVxI3w8s2dlglF9k3zEAYli
Dvz8dtgKKhmQNy15LlyRamunbdVghlSUzCknkeQZBr91jtxgLS0FU5WBAf675uCq
MGHKkh1+exyTCwcPf6ayEITIA2KYa0eSPQFP6y5UPM/wtDRvfy4diYKcNL+a1z3H
iaQhjeE2LWoL9L5zRdJd5Ed50/Ei5Dj3/zrzhYJpl+MU+FNqVdthWFJcCTiXm44V
459NmCmFVGzhBw2qo/JcXhfo2Htfs8z54flWKuu6347oWtwxg2SEfbhe6XQzmIKN
jcmITlJ6BKXbP3Os3y8ITo80jcczoGnqSwvqh5xnES+a1bPYCizj6rj2knzesvs0
9KFBI2fiTsX275JSNixE/Om2ZqVs8ge8j+tPZxTaFarL8nk92UqT/TxPmPBHmZ7D
PLnz9GfK8zn+bsiHlpDNZdCA7wgU7uugHTlVXd9ha0cYFhRjnB4OaSY2g1DypP4V
eq5FSvuaVIz2p1BnvRMg+h2wUEl6ujpUhNRgxi01qLVf0sGpXKfKtwunbm6QfoaP
Vi31UOsLZKkHUg1RbEFHUYeEsabbvS98n5CdTwwy+BWtyv6i+kqjNWJx6TsylnPm
Z/eISowMGsvmPgA1SEH0TCS2jESAdAotUzIzEonyj6Uis6UaBvTWPHWBjLqXSYU4
/NCl3kVddkpWFmK+tDv4i/PVgptu50NbiV8+oWyRjbi6AEObkncimfAiakC2gU1c
7GF7FMA47g4SM9mt+ygV6anBTJJ4LSNLJoiTezjvWc8/7dyj9dL+VK9sRiaEdQ4K
ZYjVnQzb7I8rHrROQ0ApjSa0fHVgBKH2uvuwH8Dfx57thzgPSXzXJgXuTe/KHLYC
4EQtm0rQmZv0BgCnUXCR/f54dgkVriDEqTDaGVY3RQ/kiv4Y8/Vy65UBgeREyCeW
yju0IZZcYjWDyQJGZ2fNl/3xJHLucrptyB8JeX3gzMroEen8PVZ7GALBZhpzSmbm
TZF47F14oZzI1q1alRPSUV4NeFt+YnhLPgYyml1furljlgLZYc4iGgqdPNa9EVTq
ox+/3t1eQUdtu/FsyASMEEdyqyCxtQCV9ALRmad4A5V4Naf/+6dwzH3QuQgqeWeo
FxL0VJW/x/kVKUTXABaWrlGlyFydPREcOrUfveShjw3Qc/EfUZjM6OSoUq3M/VZF
XN28ToxiwGOczVUiNYBN8eEPEow4dK2Hp4xR4gjuR7AtGA6ZUCgMee1DoA6BaF1G
lyHIWkRZCzxSVNzvKON/7hqC+Hp18cm5G+dLGqZSj9iPMMpElFBzd63XQxPbdAsx
6imyfV+KOD5XTmL4LAek7s4JREtA0friuxjwr7j0/clPXZafr6pghU5vijXmcNu0
FWQUS1KIyhLK3YyOIY9vKuhZsC1We8NW6/eWB1IrIcLwip9FgRPnpURt07Gm0ISM
Go5lWutbvTgIUlBqz386ABM0H8WMjqXged+YUmFj4A9r1hd5aWkioa6c8RrmXdcn
/PA1hfV313qYPXEG0Ij25M9sKFhdrXA4qOCfQAiLpPNC6bJGE4ye12PRYbhBqfcd
R8UEZyWasspp6d98QdNt/dbKfITbON5wm9B0xLS5vC9esn8hMJ4LrI5LRklJEKsa
ZdssyziklzFXLnJ8EoK4B+4wvmDY+IlYu56WcfZ/6TXOs3zoQMudQcDZhcXOnCEt
A323WHmRnKG2agFk95s3vSyX6bv5WNogtYenHsnoqQHpOFq0oNwiz7RhDVbJ9FWz
U2J6sgy3Dy07LQ1UWPwUF4/Z/LoMv2ZVg4VMgYUp8ehfa+BfblKKG4FNCMv9vBZW
48XZ8GKmcQwhAekIzTQiRNK5NcfdtXZaEzNGW7s1RGwX/aWGhekTmMzY2PxyUFKV
CHnWqrEo8tzh7b2mScsy/CQn/9Rd5Ug75wRbEWkU/A0wTBTbNyzd3bKrZSEXnSOF
FhfF9LKIsMm3y45ae/SzcVrtg7wSYwxg8NxDjzM7lGloSqXbJIQOuuHECo5QCEVA
9RzWElssLRsOurlaref5axZC04771UTjOxa0k1gHNlFIWxyCGcEsBztilLewMCLc
X3zRHP4HeTQG0wAUcotJl6AG0rQQLjOjQbrCqq2SvkcEAc6woMWckfrv6/5CWeYq
+6wV0MoBdl7SYx+oiKgtIRfhOrnQyD3glZz3dp0GxTBnFpnu6u6oICUMNkPS94UD
lW8lziF3TPZ5QMVCptIj5ITRrYV6FJHcK1N7A3XOmXvtUinNRFk1LuBFL5VnlfbY
+9sKN1Yb7FJNthGEsyWeEFCMuG17UoS4pbXS1ACavSybCJg3GS0DlHbl3Z9mw3+n
0zo4QA7xK3GBzt92KhUF+bx6k9cw9up1ECNlXmpGMv7uOu8BOwsDd9p9PzU22pNO
q+O4VwnfoKGglWkJb6K+YrfaWJHJLxXDV+Gv5OeO8WUtLUSXe6RYClLeMm9I6DIo
S6ciXp+qFgyByRSV64ePirgAtJ5OXEWmF2u+akGxGDB5UZ0VA7RYka0UBdx1WvIp
IREIbMZ7JWlFaTkQPRrI32cUSxXKgQ8iVBLku+rQVDS1yUOnSD7eZXxAF4Z80SjR
HsxZUimfJSQOZha1mbp3y7DzJyDejJMp2Hp/RiWAZVLEt9x4jh2BwmxG+AwXoYGH
5+WcvJvTgTST4OMtKpUxKB9sRJ92Qpkw6UwljSh5HK1dV6EpspE9yK3Gc3F0XjAI
Vw3RWHGbWvBjHwkhxPlP0xccJote4yykcUEm5XoF2CoEZzEyJ8mmMix3c/vyur2P
BRbH0s+7jw4FaQOAISO3ykeE+E1hdvbCWcs363Ns7uAIozl0dpkYJSoyQVAVWd+p
oV3I3XeOJyBFpGVMkCmfC8anipwRkQEzA4mSie93ft2x2ni5YBO2mFuONKCNo5T2
0hmwU/9YwPnmFmyY4kqNe0MU4SCAQ+T7p79DWI7Y8VAnmVwkuP9L279MRrVUXUeq
8INFDUcQ7wDE/FDNb6fjp45qZcPLSWjQCcO0UZJFtZectkgvoqd177T7zH2OZ5eN
TcZKdMUr2Sz+HRbTN13nb30eutBHmZ8QdvOFlKNvg9oSCwhiWKixEshZvzwsVqgA
9K2hoZCH3XLlAeQqOOhmlR7JkcX7Xb8MNgVBWIwrK3Ug8Xxn+tz1gb7eFt4bYoB1
rQUiL/wSmXgGIBGasDRB63XwpGRyA41pYMDA2/9e6mqxNHMusD4K+IA9ZnzQnlnW
MMCaXRt7utKozkXSpWveSFbshxEdniqOQNinGotio68yHr4JQnL35fojqgu55OuU
VSHCP+7GvogG299APov8kkILBwdkyVtk7vw/eXrsvPehza3k7hW3vKksylMOQ4MU
UKYhFdVVCAPsAWcrIV+HT1wO8Lhxpmq4hJwH2fZROT3UxX0Gl0g6ptKPBA8DQ181
Wl2p4slyiBzYCnKnaCcRI7jRBhLKoAL1arhqbQjY5DcuB/WMhF+DaeHEHK4FHm/k
O8o0L1Q8jLNICwO+tv6BzNDjhK5+DGrakgHeZyxITZCGhNOEKzWdVZT0t5Njuiw7
b7ZrCnmbhrqApXYq/bUR+L5DNrfXK8/h8Xi0nOou4brKdlV30yhQ8t4hECddf0B7
X5v2oa/34ARDki92JzZPeLyh0wfGJESkD+5Yxo7FTW/KqAjA08otlkcpMXqP2IMk
BF0vYPAInn0NrTrBb7rQkCSx2kDVxEzLVU55KoZrLfurU8fv3K2zWEAP7li0PgAR
YT4LUI7E0knW3p4Q6Ujj7SGWaUBb9PEWDF5gE0qxhFqxBdKhz+6G4m2AAwiRE50I
IRMVSlwQK3ZdiIhy9OjLLTnU4nissSWKPk0JPpy5vLcOsKAQWd/Gg4U3jkHWl5eJ
WRHR409pP9JAQOzn4P872N/QupT1MkRZvcwMScC08zd19uowu13JIwrZaSPLEtjZ
HEROa8krBOKQrF8OrckLTtxUHilVuOvZqvUAdfcYpXNYlu0ygNhDm+lwZuZsjEf+
2OIvFPhDU0RDGe/dzULEMhTlpXefjBtwgb4khzT/LARLNNOHR+Nlp7JZ5O+6LqWy
sBnVEaot0ydE9Lmf6eOmqFUit2HCppVkPJiRh2zeWakRZVEMONtyCVVOmaVipxs6
qi+Sysn8RSDeE3i33Xj8c4Wa5ny5ZqblYcKEYpg3Vdh1lQKNknNydksgImJ7k4qd
uiDgQof0k8RRYWkx+HYUspg1vztcVWU1BGkxGjzYb4dLjAZsskrVSvaOg38yLu2C
rhWrqR9zMhlq79ZixN07hKXPfsx0n2CJhUisq6YVS2NR9csE6iDR4JbTHvoEtuuy
gehnYWkehpvBZaE9plLXnVd0o20vM0kFyzmeUcTP9g+3n2WZzHifTeRzSh8Lqur3
4/CnWoO5paYDvY429iRpGoQDpKcv8NJ3tgrKXrq6u7coKq+6+hSLjJuBSumefpEW
50TVZAPG1y9hF3J8jZP/Xubo2dSbIcudKGatjob90Y5qIgiG391s6q34+Gnb/Iy3
Hi/G+XQSW3LrRKsR67NI4UqLBxhR9RVhv61Q/nBoxFZWLqgv+8+cRVTQ6JAG3zH+
e2S2jGZNgDUZCi5hWtpfdNC2M+CgHp9Tim9ESPsdtsp71ze1XeusomfQtKshRDbL
OdlYSvnYGPQBQvLTwUuwnUUGDu1RO0pdh+YtMnuYC9e9+8IMAmvjTfLMn2QiTCjt
2taYzDGCPffbskMHvE4+qsM9o+W9QogmpuxQz5Wcg3PSDdQOir7WU4X6lMg+ECaR
BnBAq9pbZxalKHWkSO8Eyncn6zSHZSo6r55JkoZHvvt9M2DgJDkXVKLKE9UFsZ20
pb57ivw/erUAM3Yipw3qUJE8thG9fRsQhmWRM0oS/s6rRuCpeaAjKptKSkzpSOET
kFx5liftMbXtaHJPxNyNWFaaTRVJq0YwbTtyHu5xzFYQTlWojpaVYVQN8CBn++SF
xiVhaAuONDc6n1Ngz+nbI45XQFyclGbKSzHUgDpVIGaaj54/f2x1SRgDMU3GAQEX
79VTOauu8jz3VP1szC4qzOiK/+5p5uXqfuUmVzfQicy13aEN2AU4ePIlsY9wrmvb
tOJY3Vn8/0GzWTveCZgW5l4AuADYNGsyaRugWJftPs+5su8vEMlh2mib22kjNR+S
cf2E6c0LlCc5JT2f30YCTCAzgcTxUUV5X8WBxGsMm2y7UEWQNrk4A+QnCEAIGg+P
oXdHbvGAUMIJS6k7JNJhgbil8RKNoKFF/HvIuFStgnAuxtDxCVkH6/JPhoFA53+O
ksjG874P5tpF0D5j+VDtXGD0h2JlEQ+yxW3HGFZOFMxld09oWrbXIIlLveAlHF80
0wKRY+no+2YODThKeo0L4d52/umsduAjRO0L5ILCNLVSu3kXx7zXZhKraogTFwv1
UuSzeEiGAGH8+jmW7US/w/3WXnjR8IizVgR9CgSR6t6OWbhZo4nqb76bWvciS7x7
DRTUOzjQgoVa3q1C0a2d93pimKXpWsNhpDKBfLYo+JgH7VZUwl7NVsi0IJoOIaIh
5ZNXG/z+r+b+9bm89IC7cGVMyYoC/nd37lIs+pXx8ZtPTMu41A6H5C29k0cE/tHL
C9jRWzr1Sta1b7bqQBxCuQiy46utaXg9ZHARhqybZGZcVDukAoq0L6UMWDn4mkrx
+//aM0u8QhJ0dwhDH1KjyLebqidAqr2J4U5ba/QIrvc=
//pragma protect end_data_block
//pragma protect digest_block
SwpNrZYnayqh0xd0CU7+F48vk5M=
//pragma protect end_digest_block
//pragma protect end_protected
