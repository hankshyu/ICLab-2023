//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
N1ccDw5vPZCBU/x4o3VWaKv5gVogkkYPpU+De8/ffHHa8iuoFoITRaM2Af5roCW7
/37NdkjTA3NdNMlvsbRQgehLn1MS3L+EkWR0oLkjHvxwWbzawlq2fIOc8Nj9yrHR
3MPsc51wib1JHz3qYPIMYHxvUXlr4cuuuOQmG/DPDfJdh2yyqQkEgVNFQPGCBUCn
DxQNENcEBG/CkqnQ75iOz3+zI4NsKTKYa0DjgrW+srn7Vecj+MIVgQJRPGcLtsQY
3DlCB+T8kRnp7WBmXumogqc0TCKt04vUbVSxv1Vg/qIixIRzrUEj1gKKM0pfAzhd
jztJVM2g4MVC9mwejg0Zkw==
//pragma protect end_key_block
//pragma protect digest_block
KaAoOmBy3pufqrxhdtOyjigmpyQ=
//pragma protect end_digest_block
//pragma protect data_block
JaEi4f+G0w3gv6OKyOq8fXnYXA2CrYDIR3xt6zF0tlW/2eaC/w/8HTygYoOcG0Z0
hjYNTaDN2UjLzYeGhPQiaHymaXvWy8DY/V0V11EDrPGztD0C46rmZZvIDqPyBU/C
AymoSWZ3/+kg26+SIBgB0H5ZrHyY9S0BkYxvb0IPYpkVYgAN4fpR9WGhR80Ml2Rr
7rVV9RsDqAoV8nd/2tL9iOU9oBdYYuN9pkDgqVeD6Ea9411txp9yJ8loM0a80+bc
pFrmyYVqfpFsA5v6icPQv37HUb8UjKoGMUWl6XVS29u5Mfb8bVlfnROjyYc/5fKl
tts6dqvVlah9J8c7aZVp5us6nHubIAJ8JtiB3moPUld72GwQ+9bn+3CObVagJ27j
KoOICGdFUfm0MvQIJluCQENip9+R2OCPKEXafA7MoiIMVOqVf5R1J4y/w8SJTqR4
cN6RTB+5coQW6B0XZgcYZZrupIQLnUwM4R2k+0qkbEcEeqQArx9wZ9AT2sxlTe3n
ODg15D9tGw40NJF2aajuH/od0JUjrD0ZlYtAhNkn1zpiknOTdM0Z2gJU25nnCn1+
nOs1P0YPEHz7xwD3UFm4IoDYT5pZGiUN532IyNKp+XE72M70v1bSVX187FgvKW7w
UdxzH+0VxZjL4Q/AlUh3UrNKt/aObzkFVspxj2Y48gRN5gDpT9ae6Avud8lPscoK
BsbACUr8AREFM8mhdI5EXdz743Af5glPD3la4/VO7uPk3hnaFKbjh2/H1RCPZTCo
KXxY8qkMgikxV5Q+bhuIndlW0eeRCwQLYRsusBKOorRZw1gwtdUGV36qmR/46/qU
+a4kcgMB0XkrIQZj7oRWwrNTth36Zgpvuwtcp7JKqnEpr+8PYqt0NiRaZZ5nL4PM
s905cCfMjsLnBy4b0YUkD4OFrPIujEtzdxoOMBUCP0amPKjIY1Ga4E9mwP7FCig5
wFBVYdA6/XCIIzsdCvYpy5LHmJZmMEBxC50nz2TA4+grsMYcGkTzK4CWSiytH0ee
pyERd6aqdRAmXZVgZ8yLJ+TP0fflKUCZA9lZTGLWrpjJKwSmHuzh3fdOf4on/Akv
bB9AVPwNLBVJVR0ciiQ9xjEWS5OuQ4gmksdF4ha2MNqlmVLT7kYWFg1pC2jyBlPC
Y5MmtU6GNZ1Q2nN7n3oziHm2w8CaZoDcUGQGAf68AusROimbAIiPZnOSWWyrWvmF
w0dRU5h25CrBu7whvrjm5fxfNvnlXuXwO+vyRVJavRdfPL7sJI3330iQbqmSZMsW
hDI8p4I/RD4aR6gHVQBd8tK8+Siik0jvm4+P8Pm22G9AEGFJuiMyGF3Oiuactxgt
Mc1vwREek5JEr0Q5+3VK0f2RWovqfi206sgCbKFSm8pRU64X0Ly2RHzf2G/uO5Z3
WjxAm7p3v61zUTuy3/UILDc3J1v16YZnhhTu6YC1XHE=
//pragma protect end_data_block
//pragma protect digest_block
BwuvgqKudPWNHr5BHgilD7/d04k=
//pragma protect end_digest_block
//pragma protect end_protected
`include "../00_TESTBED/pseudo_DRAM.sv"
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
ZxMJXU3M9nYTNGY5Xk+rtx3IYyqFtvSL4nVzBs+xSfrErMigria7H+0/NqNqvvs5
aPYj3SDPuhFtSapg+GZUDAHTYJqMbt7c44RSQ/rkd9cwpuP7AHx83wayUUv0LHf3
mPuRwD62vcgEKWV0uw+sSJOjS3/QL6FGv7klj4Tu00qd7pev5Rygt9r9pmLot24n
C6cHeW1NIDXzt/wAQn8RcwZjNajRAfLzAO/tXiOVhMV4mzqDdxyzlPHffn2T3g+G
/x1j4wnHGH5E4u9E38dBlO/svoYR1dcEF1/pPMbNqcJtpBldqPHBav4m9ElNTroV
srT+JIP/0lWW3DloRqgOiw==
//pragma protect end_key_block
//pragma protect digest_block
QllXsLOiGl30pddQtOr6mroYRdg=
//pragma protect end_digest_block
//pragma protect data_block
NZJWUitKDLi5OFhgLnMFhoDQl3I0G3jaUYNXEXw8+LE4ipwVTJ7ED59CFAVLONhB
W7by7jsdX/SbI6l/nGz8tv91c+b7O9U44P92lLYx7lBudPhWhrQx0pbOcrjDPvaL
T2W2H6VXYJapSkWMGHrfXOR5QQKorkVpR5NUnURRE4WEl7fO6emlIjnTJK6/JE0b
iDj2Qg5PPDK7NP/6nbF+As2gV0WGPFmrD+JathjtzcIe0OXIrWAx8ija5Y4PdzAd
oLkXFlk9UyTfjcsCaG1aIHDWm1yDH9Z0BWwVPWC1CgnHP1YgV1BuiilBEa1K1SIF
e3E79BJ/K7TDJiHRUYPG0Q==
//pragma protect end_data_block
//pragma protect digest_block
x4n1npZZ1uXgMJbbu7S6kh+KC/M=
//pragma protect end_digest_block
//pragma protect end_protected
`include "Usertype_OS.sv"
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
aD6PwsLuF9lmAAOkweRBV5RKR8sWTg+lQbLtEvfl9P56sJncGAISCI5mMVKvmPxn
Ld6EHoMlKJwZJ+WvMhHqrfnuYBfxcs9RM2MLM6YiKXRaB/q3P+ZBf5pdPsqtCHTO
hw1EBQT+NrqTPjNro4ztByXpuuvpebjK4k4X6Z26ZDQpJBwu73hNNktmQA8y0b0y
mUd6xLOLLZxLZBjpy0wslbKjvhoTMjPczmxcRSNuPsmfZ8+vD3edUDwEQhz5ujRB
3qZkgfSZ4R6i2BDxd0E6NWRg3KJGmd0IqvrV79esp5goH44N5B2iyRKwVGFcNAW4
TtqUxMcWqqoP37s0eSTw4A==
//pragma protect end_key_block
//pragma protect digest_block
MfZdbMK6+DLn7isx/uWASA3Nit4=
//pragma protect end_digest_block
//pragma protect data_block
yDaK/4uBSz3HSt6uKkAXYP6YqV770+wrpfpceLmItnDexpSsmPYaxR3TX2jztcjV
K6xPX6REuC2a7YHGuOESzR6ubeAgJzMN6z5pNPqgNiaJEIpmTrYPEMC6iICJWQt9
g7N/Xe/Isr32Lq5RzsxTjjnA3JrAFP/TFr+9dz066ObSapNvgXy5ngR0/iPmv4BV
B8VHphJTsXvQogpnDNy5YhehkRqwCXokBMWayS/LtHvGcQyjLa9xF6uYuTZpHLkj
xdl996cj2n/q1vym4FGk0Q9Y/Q0AfETzBd5ZXZy7/h2hxA72UFXhOs2qMPwfiO/4
tJK/fDJElUBpCe3h0XQxBFEwTJCEmU6Uze45ZnYJoO5L/tqO7Fnwz18xtdDRyNiG
P9cPyEPX4nv2nutAqSuflQ2GUdYHazWgoUdGWKr0wbmmCXb6kQolgrRUUpnoPCz3
+K+EBCssvj/M8k1HmLAicMuJP8UttuDeb+vUJx4Dc2wO337N0zzU7Ynya9/Bmm9o
C17N+V60qdoaZBGfZ9VVziWuOdkU/YnS7aIp8axEH0scAh597vN20W71kmq4b71/
llFjp/GIbuM7efPLJ9JLPCxHK6JLOCY8IrvlKtqnj8dG5pnPcxoJ/qT6CsWPm11Z
cEmhoHaEuWMsF7wHnyJj1Pl3+MNbhr7sUINN7NP5CkJ1+WTlIdkM36u3g2M+Xo/c
0Ice04lZC782fBd1I1XZMv4aW01xRiT7JLo4+EJVEKrfZceydN3sydm/IG+pnzJd
qR6NLgmRYlHkrkEkSAKeWjAblT6ZJj1rSwIE/jMoWN++IlMEy7to1cMq0Q7D/t3F
kBp7tR1jZK96FoOc6TaUSQ+OIMU1uzJPMlrKHe9lJkhJK969G9n11oube6kCrJ9B
SoSjIRn6nnikCt16/xg8fP1l/mTx8y23yObNqm/+ymFkka2jbnHfUX68+J1mtGZy
PUuboYe5IZZhjQbUrcGgcaGYULPe0HZF5PzpQRwtNVzo2PTNaCb4b5fj6DiSPAQB
IiN993q2HqZ32wBx59Pe+fJuIMkMjlMsfTem4UYLVxHZGZe9TKv02u5WkwncZSWN
M8/v467H1dm4HrwQn3DIULY8/KO/x8t/Zv783M8Jha26QBR1EkCEOsfl7L3mkzez
5GGf0gm9BPrSY8ajOt9S2DBcFCKQexvEYVAeb0GPg4bsGp1BdHc4FpXoiNNYevnp
CXPRb1XLxnUB6GjCnbvyDOXSUBcvnaQ2Ji9vMmKz4/e68G50sq+4e/3goFxQBn5m
YNyxAhqfCT/FxdTWeTUAgefUCpElfEa1nNUIQoSqWi5x/MgIFuU1zov3RQ0kyegJ
MoTLg9kMonM6T54oZ+KVahaeNVP4sY8w/JZJDqBCIr7t5Wqum87xlCL00mKDiVd2
ZvpkwozwCOVSBucon45f8GIND7BQJDMxJr2TgHs3aUy3Z4RtFddVg8ImNW4Nxc1N
p1+/jQX23nUbnkqIvzYjEuRhJY6EGnL+GnRMfca6BxwhSMFj4uZ/YAzv5mm6HU5I
6EzA2/nB37hRFyZ2fSXl8kKDDrBGgxPxC0zr//W8dGh0xOx4B8+b5fhq0MenA3MY
/2rkJThFX/6CxdouSextq9EqnXoWPrheFDlW2DQVs5DRncJjj6zEqlioz5ierU9z
Cm10H+8k8RvpLsxbT38dtEDtwIWbe9wYamPbzhtEsNAZg8f3MeurlXHfm1aqG7zY
Pr7USXQmphNLfAc4mjj8kthXKO0bAqMdGhuoYZsfi67cfr8pPhc28625QpCrGWtP
sO1SRD+N7L5OgHoTKEAk9DsYSFaWEQZNrPd0iDnUALuqdwXqQta2PysbFg/D3mHD
qGY0o/LNGhNONwrYz/FxyaK7u4O4JTEbFH4BoI4GIKjFmXnP5uKu3P0tNECoV242
spj/V4ZuyRZorkRVztdb4OADTTeKGQezEcLAebvtPUFFoArdafwDa71TL/tfiz8Y
/kbYVyKN+QhIQplEDOpx+leC3dS4h10O+34Xp7s8ZmSSDTP5yu90Y/SrZB4lPXGx
AYupT5Jbljf9h6HCwW9KyBABytbv2lIffmuza5BU1xMup73Bfyf4XCR9zPKQlSaG
X9cw0mYv+f2GjN9jA5nrKiUmOv3CLozQKm11R3GWagAbJbzzoU+D9hHdKWsRt2F+
ju19VZEonI5hfwyR/hRBQaM36Fj7gL+15ehVLuNVRgJx3D88GBhUhIDhPe5WSlwQ
zfnGYkBGps/6kJHkZH5nPYp25HnttI1aVXzVp2uAfWdrBsIjYvOxJQBwLJOAl1pw
XfFB1tLkgGiTjexuvHPhMplLpLAhPSXmLu9oNGe40sY5GJNhL8un/pXkA87CfguF
eAghUnkhhNq9LZQwA+KEMPqepBa6ZYGPkfsuQFE9F7eccwG3de7Rky9t9yTjN0p/
XWbThsUljSB931NB7VePfqOqlH+bn7d3H+3VOE2T69fczBn7/sxgXL30L3egSsB9
muf4TbiJehasNLsSVhe92d78PmwP9zlCv61C6b4TOyHIUifdDHPSks8VBZebTfws
MVMb9Twjngl1zAuRTi8Moos6zWDPn0d5GlfFIk5PlFS8BzCH8UUg/WMig4G1iRoR
F7MuUGWT1UEcr32QTbIwYbFB6E/VJ/1crl/EkFpJrFnWIxIW1wRS9G8Nn+IgzvXZ
m+LdcDYmQk5gvJaFjOyt2W8bzcA0sO/qaqoolBRrWAGFW5clWlygBmPTekAI6xRW
MQxuoVbb6wvXj0bg9/rIgsCrzCY35l+SJXXrNbEf2s6oZ7eaqoY9spBlDKwlWfaf
shQvl/g8H6GW5otsLh2U75d2GIMxM+BYD0EXs3WEaQuYrB/8MPh40eMzAkXUsfYh
ycXJqsrlyhu3Wm5cNS3pj/MfbEYftESHWazCh1dn9EhhKRMSAdbgKgSS7Zm1wSSP
rNi5UeEChiGPPgdyynLVUGbQV33V8JyDSi97v3N4rRzFyX6upXU52ApCKmfgLySz
O5NLYOb0f9NszSLPOsh1uHV5tgGwjzbLVbBOOoGcV/NRmDAV2js5XM6zYjwkxyew
tHQto5LGF0aoIgo3v+a/Xep1CxY+KXoAeX/jb1EH/aWLe8bFdNx00aSUXUookrl0
spvY12cnRHhJljfQ98K87dnhW/Uo9H/47AV8lOHsUU3flTCGUaUdqeEe+VnACJ2L
pWeUGwjDLZVNUslJRM26kqIqL3XufSztdm0BkkWbSsA1YYSBrlTFGXpIs+u3bGjV
oqxbciIurKOe5+C9hX3Tv8fcT/dWtKOt64vDH/i7j9PWZmQM+DsAl5KIIKEAac97
QQipMiA4/mAJkTuCYBiYfFMmdvRCRC68nWWDrt0EDGRmEZmvfWh/fOILLT81qbPp
psIDnXHkMylGyt69m/5Ch66paZVwkHdQ/p2xps9Y7WQIQeWj48E5NOQeL4mqao3F
U9ObTkzU1aulausFhX5+9cggxUVFiF3iUUJ4ixK22ynWppue4hNRpHJUaVIK62YO
DyRKB/4uG7HzDTPrDvO9Eue1rGzPf+n5Xy12q0E+rbU7i8KJIrnJJ8Txg3/9QlX0
DhVBh8wJmuqbls7CggOIxKFYSrr4ddCvqY6OOTNVeKdrMR4ej7mRfE84mZWRrXqc
3+beyid1Pfhp6tnM3T8zAf9sexzhPIEG7GJ6U6gBIacsSRsLqI+Bx1qAat8YypZ8
sn2PN3sZIpf8rECNFm1y1TaYbQ7m7mSy9HlbJVe2F0KKfcr4yF7sURx6LpKZVoTs
OYz5CwjTlecs8zKUmYGNDg60dnbMA72lClO3MhM+sD33wVBOiObixhO78bb9un06
hR9i/ke7tguEYCjj/77lmwm0eabErY4718wOLZhReCQMzjLB+1J9DtvRBDV6QOtB
/haeZxpsZG2J5hYu71diOYWZXPqKHU8INKoJW1XE61k5onKY6snqtkb2Wx+ouBbu
cji4mjNuAJ7V/XeGJ0fos/KXf2YKbcx8yAX2hxCYroX4MW3Xeug3jvEU6wy42w4y
INtmRP4ox6nkGGbz7cyKonizjReRjkwN4kY551j+6dXrZoJjAMwdOM3I4jrc1hyu
PTKMRYXr6WgDCXkmBP19Urfs7x5qZvk2Fvw5pwm1IhYCO9OWIlcdqzwlaNnb2VgI
4c44J1Ypnv56F6nhAR02MSq7qrYyFERcZViiXyMab7qCkM/m5sPE4N3ssc7MuDwV
eOhSSd/1jtiVnCfBp9Ge/tug6tTwrr2QgkEyK59KVMjbCzyUc7fFve31wCZmESQC
wxy4ImlQZC78l1m+G0VDRGp5uMqJpdLrzwOTe935fmALsYBrjTP+KlWeZzEIrbiX
Q0TsEAVSoa8CnvekR8lqqj53eO0+/O674eFP9Of0FEOskJy9hxi186UtQFIvNbiE
3kFHTBvotfRrel9+xo6PUovuv9x3clspjmkK7PUCXrLDt9S0wBrYnItrdKPuTpdq
6pUDV7To3Ugrn1FczeWaNJZHk3BWDjOZFRCZOKUVCw5nCNS5slvM9HaH/hSzGbIr
s37msyz0NM82AaRVU4YjU3cXipoLHqew5sYZMnREA8g/NsBUfPguKWH3wHDngQFr
dXKCYkyRIyppwTNqD3csgvbWJsl0O6JvXCQ0iUhm0+SCzoay9juFRUjCdTkkMtR0
wes7Q1VzBuWKlceVlmoK7i++P9QWCSvoPl8/eLggqm2EKzMUWdbMHzVDUc8Yy8tx
Q5sBnq8Nw5cgDSEa+yZnlFM1ScYs1vd1h+gOqOrLBEaKDgrsjakTJ0KS4zk7YDFB
ZYJ/algNuGVUVdf4nwBFyq3pJHDW/vom4JdS9bTMUsEslshnF0d/XL9YH7QrTSWS
t0LIWY2u/Gig+FlCKR62Eh2s0ZUlsonteydBa9A7jwagdDPKxtd8lO0M7e2RGgiY
dsOcozKAhHJrBuwoUdirXORGubxdg4dPGWlm3y78JBF8urCq6ZhSJs4KyUxp5O5i
aN7CB4YczZav7mNJQhOvThbNIlWrNlY4/o5rZ+/hg9CyALCeMYa+91gTxUq7tTKT
nXSJk+rzWLoYvTJ//F8hXfiDvJuck7EL7Eq2C+4nq8I/fnfsTxYZnesJ453md+3s
ytDpE4vBUNbM2c9bSC4cqRryiSwnrLAPhuJtZs00huMe4717gJ2eOTs+nhcLkoqr
pRhZY7zBInQ9AcCTgVO6DbqxS3D/Rk6TxxTfD6LU0Bnb4XSKG0qW00nYQ76Si2RZ
HC6pbMH74qsQunhuBgybKFtbrFnurEa5iaK7yIp4EGzUc6HMBfPwbc0GrRO1WSIl
1t7Q842FHhx4qJNGk4f1Zu0UBdWhbqT36WvN9ZUcT509zvh9+AVGLAhW1V6Xt5Px
h4zGRPmkdwVVgf3UiSGau6XMYsEkWw2MC49FB5M3P/9QHM8Z3JooF88ItYu79mpz
zwKHWaMOyFbOx3Tiw0ASj9DogOThxE9/tSYv6RVyU1DTJ83AaE5lKDH/vwlRFULb
PWX9SY2eECvmkhRc6LBgUvQmDqVdidSguMtp840YSksfGJpsT94czkD7EnLe6dqW
aqIusSwkHAMj6GgVtwvGVD5OAkogAts7u9ZN5j7iXsNjnf7RUh5FWEsnJT0oJ9qX
h9OR0DAO3vI/L8DfEIQ6rx5JnjqzgXSwoudnKQ05+lnkkcXgAErrvQrf0Y5Z9ykM
9SJombMN8gCbQ72VbMaNHib69ap3B8X8VbRHIulY6aP1+V8CU/cF8EUubD1oqYhZ
+MByuReI0WPDPWJtGn22jyZqhzyUUqLXhUu40ZrFs+wyFDndIPnGEMPkRup/z7z0
RKX3wxxbN3A9n4tQmSXtV6UUetC1u6R9UaP/JUSGXi9p2bLVCZ4fAF+qyPZEkp5H
EpU+V6/16VTYXgIepTsX0TBtcSBUbzrjZhrCdDf2CciIyc+a9+ponSGzFlwXly19
Bf/yMTyYvCj/Z5gckB5vo/33H816KcHIz7znCzhSKNqyP2aWOXuLtM5VOjifjB5x
k/+oI6c9Cp0xRbDAVfV846q8bvtSG4IIkVyip0TX1NV8jqzhQQTedBffIcbqb5Xd
cUeTCiqVb+p3HEE9lwmt1khqHWR9d3d9fngmTY22k4fYiORr/Ba0VDAxWj3EarLi
1U3Lmn5QFFtmzmlk1G4yROE+TVObGWvOrJzjlmgV7XJRCbbpi460lr6D96cRPckn
EuDzIVP8vXWv7Q4R11MT9ZbXRvMMXwTuha871Cw80Emq+Aol53wV/GhSLG1T7OhY
0xSk4wMeLYL0pccw+meJc9EzodJFponPm7bMbZMJcIacnvdAlt6zkmaMjmVJB2C3
NvCUy1bU7MHApt1ni+R6cqdX7ifLzhHpRdfWzgV5kMsFZqUkUODVONM/jX8xrZ3O
8IdDKrJ/+HtyvEjm5Hz1/lGc7Dyn0KwTdC5zgtPXUb2Fv84AW2/tNfzkZdXAwTNR
5Rimtzd8xTSzN12mj8kZDEVfKuauc+d87JGlRC9slLaHC51Sf9az+VHC3AwzmAYV
A36bD2Xa/VOObp/5uLbSE0igbY/K62iANWVXNY2iOZfZn4cqe+sxFnxkivXr3nv5
BISK9mBIRHIyvWIxhZl5oBKnflcW7AnjVaWDdXnzIpQNp3i6dbpYUiW5/xd3tFl2
2fWqA8AA3Bm+WCLmt1DGNFtD4X2d9rnVYUld+7AI2amNzgcAwKxN36DVr3ws6/pN
BBpcIRfyqLFQuX/gO+O9rDvRKX+sOe/JgkCdHycJPDXYOOUD+B42LRqiIE8ls3eU
W9rrg0/GTuen5+rlkpecgbt6miQcObVkjg4/zeaPw8lKhLuvYcpfkiso1tPW7oW2
bPXC/Pr4fbXRp5eHWtxdbXREgPkGjqwVohmwGh3uRq4l4JwhkBooxUfIbzTQnaOy
JmNwaVlX64LhAcGUbpi44NCJtt2eJR3f5F0Axr4zvkx6iYsHNmoRr0U3h5lJiPha
K58PCYxCFwpRzY9WGoCcG/g++1GJvRWGU1h2Jbo2/5qQlMxBNmymAf4g+UVKV1WD
eG1mrumT9BN2ohs5SNaFFSmsOADJB4HxCM+t04YmLeInbN7tN3jGN8Y4RDYfuM9P
c1ltUqLtqpGUu6i/X1I0NAKdHuvFVhWFLOrBuV9eFIv6qs6fh1U1bZWmUr1TjHfP
zMQHMBzRbdl6e1kN79hLc3M1/WaJTSk5F0ONO7ejo4b0DQEbiJCzGa54oNJMDV94
lh6weIZCsZTC3tYXpzC9PC3oMj7FMzj6KyWudRFFHAkmdTyxPbFmxVWM6q45Xs0C
ot9QSdFM1d40N2WX7RM4TKXIw2p98XCo8OqzesgJ30WkxYWYKf8Yor7YZFji6jUN
SjblDXdA8vs30WSS61hCBwzt2LTTyhWrbjEBFmWy9m+l23ipgL1z/NTGK5+GDwkc
8wlxd5kfic7pZ5/+29yNDnidY8I6+ru/zgBNJtRPZSWLZjTShnhjPpM21VDdZqVt
QwLy26LcU1QgQ272MeNGW2QJu/IV0YHdNik/w0jaX/6YJ/CWNI9AVO0UfY5Sz8gV
uerNXPIAiSltNNS2BXlmht0rB0R8SGq1ok/KzqSYGsgtvwiWm1sblZxgEZ2tUrmq
w0icskHmPZY1E4LyXan4wTk2tDLYPxAqu3EmtblKCoc6H2Pyl2zTSlkR8kmT7XJX
Kgu+nEhlvjeHxFgMWWwvK/CpMXGF1Gt2lpYYLdIgF3jXDjughJZgmY9kdJ6eRZY/
KUZhLQLF3HyTOB1Gd++8b4y3r7eYE8hJ1bKADm1eeFl0qy3hUN0jEHjaLcs6C5h9
Kdq9w2MWNE/i9WK4987m3GUa/p3gx0ozmu8dU2s332//I1W1w84d1rNwWWKIlyY5
t+tIQMX/9PrtZUD7ZU7tGby0ktJLskBQ3pyW0i4koUTNOOVJUIGK+57eQwB3CFei
T72L5lRLZ371hykbQmxHu3JLFfFHLZV6/AIKHt7Kg8Lg+uGInudsqyM24sSNXVZE
bFRG04IPBr/jVM/w26Xvom2AG6Aq/cAj2FelueZYREY+FCU+I9uHGdLdKTVcebPT
rY4n7DIIFoN4hsc+IF597IOWMSC0vi4xW6DYsV3SlrpAaCKshkb1lcACXO5YGAuB
5wVamI3WBgoo2gjbrVe1AXm8Lf/Xo1xACQ/EEMcpS6h6dnqxm6Cg71vynhipR7uB
6tthbtQ39nilTBM6ByZHxlxoLKplIbct1RDRoHdMPPF5KcgQxWQGGSkebNH/ajjT
EJCgMQl7n8l9D3GOwuS1rhOxzSNxpUszTJYQ4ZVPAkLREldUIPKePdpbNb0CAAjT
ltMgs3l2uWGDNpOkR2PANxRxDiPDF1X4UuaClIWaid8Ss1XEHgPI9RXe5R1rPkDp
ZuSy8F7hfgJ8vlh9G2QVCFX3U/4kkRtiVGpQ3R/5bPzXAtWOEvqegnpB/NJuVnzD
Iti0GeLMGBj/VEl1sO6iSLthfWwEXraumt4EEGM9ht8o228yy1idmO9ii8kQVRBx
sAqRgQqt5UfD9HXt8mTLkfeAVxOrZ8eCTUbUVv5zaSPpzw8B9Ro9uilHqNY8Zr70
BWzoWtlaKHvS7qt1HjUWIqdTkY0gbh/BFI1aHvFvB9aQ2cWHYi8jjkBXeLHq9bUo
+x9WRDhYcKqf4aF/fMs6pBbqG4htUhOMp1DPO1S4LNga2hOmrA52eEqFU7eepuiI
PQJqkv/qwWqe59WI5dHlRowufOw/X6urO7KHoTqqU3vSlSa1Lypv3QD8LshH2zIu
mmfcJ2qMrTCmOApIHqc/K2LvV3oqItc0Y0tosv0NI380TpzcuYQkEPxvCY9VaH1I
ZLN3sapcMj4+5CmTCywETV6IYW5xjqxjGGVzHAJhFCo20E3zz3fobxwjlEnAFqYD
k98rlJiac5dLzAssX1tm3m9RLIrqdvWw7RFtZj+x13loGbKm5dqan8Q2dnqL7N68
72zXzY4nbBkrP5ylxQsBuSWSEMvnlAr+rRapk0rinaMLqaGlDi8xsXi3oPbFREVu
7nNaO8itYs/6VWkt7vD8vFobaYmbP7ejWa2zXJxkmwzrudjVqoDzDXCoCJibihd9
O8+Et+3vnZkm7RALvRC6r2EY2xydbbJuJj0o8a3v1kv3ne8j437Ch6Tx0d25dbbc
S7jF1WqghfTGHTYJUCtY3ScubEukg74dSWE+dj98TQH0YUDhVYPVG5rprtgAl660
maJcyCTVzV19MO/VpSsPU0/9YSmfZLeOaE3kfJP4u8FqYN+2f3ED6CU0wg6tJgH3
4klkRh7qcAzMhMb/DVFr/hkJEPMmWbv4bwFJ9yr5/yoXxY5eJlCDGuCUANwBSuNF
VfJgTymEM/4QY1R2ZW17t2CKKJqyHvjLtbJTNkI4Qa7gVeboBqwDbThlEZ7TkU0t
Ul3d9LpmHIO4Odye2zl+kUyaRkxmhODD9iX3XhaU2uvRVSwNaE24zgkYZt+Xv0AG
G+oWxeujcVR0n/UqE8e4Z1ICZQRojwlaiFjEwkqNETl5gpmi5LPQCI69fBjlAK4e
h2xVIRgYmbjzfNr5gjat/IJijTK2szD5YptJnlzEbzB6XYOlYr7ru/bjftAEqjtp
DioPzEBa9ZBoJusB4yMv4NYW65y6nM+7sL8RLUqghxAO88XWmwrc6jOZGEueiTqt
ZxuBlFApD5eXEr4xrJb3i78H/Aa8gBG7CJ4S2Ius3AU74M5xduZbkRK3+DvlUQQV
FXqVrlC1r3FK8bOvQF+AK6ip3o8uTHvh1geoq5ENbQvrr26yeZCbPPH30jGSVWqs
o9gGYQ33++OcQhgDCQKLO9r2BAbM/El9o3Co89z5mI1a6y1up/6TZ/UfWhL4w1Ez
xelXGmNt4tcTE1aAQPNF7fjv2Y+LVAafa0/Hw8CJ0J0XnhftkiuXq9Q6Y2HBZpax
4YI/uxbTqUuDYpbesxxk7qinFL6ZligBkoHrrV3TG7X8BGUyJot7SyBjHnISjP3N
vnKDmlaJY+BOvq+lFArsGZLUFxIksrs850HYEp3xCGkWD6oozAGMnNlLWzHhGbUg
9YjH1GC7euw50vzSb96u+4UErmL77C8eDcouUwyzwCJ07rtCnrqDMAO1QOEcbAhq
GLuA475yexCYO8nuYJgYU//pAjBYzAdc2ckM+G9eKT8H40PI2Kb4OlusKDDcB659
NNnt8V01FAH3rMpJl4OKTn+lk2A4OBkAj170OJWEpYQGZG/nAU6ZNm/0TFFBxkQh
nMa71QhdRuHOBstoeFfmvT+WQNau/TolooHhcOriSKFIO0e0qHe1pc53zQr+ZuBm
nCEAWDH4hmMM78II+Sh5SQeNL2iTKIaQXjWVVTlFo7z0/wRIOIe6FwusJDcY5E38
DhKvcFeVspcYx1pBJW5ZbYGnHxHz9LBai8Jgi538u0/oJSPTd2ViqmNPvATXkpyD
32wBzfE7m7HZXB8t5JJhnQyz5/vY9dPRM908DtkLqMRAVwo7fjh5f1mWLI61pr9A
C4mIKPcy7y1W+QQn0VlgRiffHlsGl6Jjdirequi6FGn7PFieIxIx2V+9fWb8c7xs
rnMdl/sLAq42+DBTRMdpMbWkZuU4PwjUNc581iatFrZnK1krt93XXxDNncNvhTfP
ZBgB3cJPHT8TSLMidkwutRaVkR8PC/5JTfpdJs9INrTuI2ei3jHx521s2M0dJ9do
rPTO4OIIc1pNR02+27HnVSDOexb9lSgLLJw7GKDR2ZFbr3j0jvquPNz4/LHaI6zS
tUneG6nS0c7K914EHX8plHWmN9nxyHZlb+1gavCBc9t8zd/2C+sF3ZMkoLFGmnuD
7Cdm5/7qTnxR9LA0BEpDvVx/BBVxtWfyhx1cd/kuJ0Uncqwc4M29pfiLHgOAug5X
1T8Bgc+VF6UEEsWxQdzV+EbnL7SKK5+DtsEbqMjznFqfYq+OPZCkbctT7Gar06AX
JDL8wWZETEISX8mZ5pNUN141zZZ81ke5ujNqC0vERV8teuWZl1Yk8/vc1IdfFmpZ
gxubs62g1HlNMbyZhJqUMIS3JrG0bs8E15PXn5F/7FDhLpOXwjtIBAdaEA0c8/5C
DNdcpZMABRzPwQEPSgDmBiT2GBuYwftM/G70T/UF4/cTdd6V9Qw4XY69GIK4ON3+
FZrqk8XItMeZUlYHzVGNu+79tpkh4BzrEtjASv/A5HbU4EkgmuI6KmoqKsrei3ZB
AZraTf6aMtLUsuEzh30gYNK7aOBLrEyVtYyIlc4/UDZKzAty4WCvhu2pZ4Wuh89I
I+BeTSb+foEVovIE9Pvopw2juAo2/3sNBKb3KKqkqMZuuVrl3WbPAUYlA7E2GKoP
N+DDQxEsLVz70xuBWJ1n4gDDeTr+jYB5JNpp8UEuNgXht3Q6EKq++nGlGHfQN2Lj
fHoQXbPmu3ePZFKtOXSsNMYxlnT9tq1kRI9FLJVUJqnqKJp6R/AzZoWFTBKYI/Lg
737s0elRh4fa+yU6wl0vpDoCE6FAkbV1Wv+hhamAP1FQDPt3ALTJiJxibLed0/Vm
mZyTntJGEFhVSjXsBC8Vupeg76E+kHHB9aV/fSdhDKjN+Pw3GUtIUA4yoU92g4sj
2agKNucVZosnc7ip9JkVFL8tl/8UC2jISd5ojrH3eaShyM6mF7HUsQQaal3oivyK
XLRGrPNGNnGYEkrBmMeZFDgV9MymQ4O9nXTPTN/sUylIQGwW61T1Kw/fIMb0+C5k
YHSR37Y/WRhj6m3pfYZEke68D4JEfwvJ6b34c1E+Kp2K0nIuvPNHeIT3VuLf/zFE
42eHHDlLu6ARdIC/KNodrLcfckHP07284qOIb3TtUjH3++Bkpjjeaai7jgPIg7Z5
VNrrc5mZ4Jt6hbhCqrMJCuEsK8QpMGXbb1COQtUEJmT0DYbjBioMPng0wrO4ART1
WVFuc1pE88Cd6EnAuUYRWBjonji2ifNUv/CmTmTZo+S6RK/kgZMb9Zs/8PB3XnJq
7ZL8K2BjanvXl6LWH+ahCk0+001Svay3M+a5x6Mr4DujeVVN+VUjSdPZE9l4wNjw
NNzPSbXUzG370WyzJaLtmVL+zDvpCcKWYir37y3/xtLtvf0M9pwNufr/N5tgrdmy
1n6Tr/DyyYA7u5+A0WzFvE7sSCX1xOJPRZ4PRCwN1T+9p6sGtxtWXsUivGSjwHt3
Al01YVqFkZzn/yQHCq+1mDbGITayE55zRHQayWUxdbTBUyH2ts0GffcTF1cEELEQ
xX1czSjZvGk34Ek3SIdEF6AyiPZldHhmby5ew+/ChCW29fm/ardMPlgpehWN0zCW
t3E1xWzcVcA8kIOC81W3C4WawKssGQ1Dzh0rWS+07vpc4zkdva6sdk3gphGfdfj2
BQn8nSZRHv3RU52vxrniqqxIVYsBtxLuasLs2J3yu9oRsH1pZ0DCIdkhSliutVTw
JGSOaWeLFBMGjEasq7Yam21J33z4jKldydkvJYI1hNpJ3RTioz8W1BV/fp25wWno
LqAhY4ZA+LDbFRJ1/H73WBKinBdly8Xp5HpgFjJUQJgiz+/TogaJAw9fUaUniu+r
7YA/TTSQh9+nxq15b+PYELM2YT/05V8f+dl1Yjm79cbd+tE1kSZAXUSINSNC5V10
waMPVhJqqGQslkedy734cNuHItK0hgM5mJUlmwXa+vwkjIxziWxE2BLICoFwgUPl
yBO6uhvtdPWBdEUc7QayY9JXNyHprzq/KVW7Qstb2j1IkVBwWfBsGpqj/ZPbXMgk
z2XWe0ehGXls73fVcvjFHCDwqynnmB70gQ70oOInuRkI2qW/NYiA/eYw6wVj7cbG
8Q0OxJl3TOsnr3P+qq/8c+PSJXDaGsCNMdsrQ/j/rbsH96aQH1Vj2VaJ3lvETfp1
rZkEhcAC2EcVMtfVoQZrsuNLbfsvHRxN2zGEvoh1UHbsyiWtZ+kHOj46aWRc8/an
1l9chDxO9cjunoD8F8Gnm+emS+1S9IO1pcfPMUiLMHeKjcywDAmIS2/zM1Gmu2Zu
Oule0QhKvdgqFh5333nyKWSWkSJp/h5m/jr/C6z9FL4Q7x78oxwIhV12jNj4tUY0
v+Ux2riFp7cX1frDRZ9abk/2EGqagBsgKH820UMUlnHwmoAPFscVS0l0+R63OVk8
MbV1iv0361RnbLM+YKWFzBdp7vJLmpEPkgC1+m8ZWddKRIPRi0axlFspuKerbopY
Hy7wsK7G1RO3gLLHqAbpMmy97uQLfEhttKe8/khYzBc1wfARYQpWi4yTVtQUvZ8P
/dOkqGBVkQMXfNtcI8NLlNhBPyz6Wy5zh1KbNNQ1EinjkeZGEYFMy7wgx+2w/meS
+B8XlKqAcR0pfTLzx6ADBfX6KOxJgE0LnuhxuWkSJgMhpiuq+Tn7B6A6iFfhJXdD
qzPvmV3VvloxW3beri2Jxt3Oco6joRWDFnRW+cRVFstJqnrPfUZ0DmDYD9UPpmPc
agC+KgeYTSxkf2toaZ9xBcvFbJUD0/mdVKoxWeb1pbyQFBvxrzK/NYWPFWL3NnqN
N1z9qpHAjhh/5GBYbbykD7dvKtIl7rbXYFhXxHEuvtv/Mo79XwpoU/2vVMPeZ8cJ
r+BZvtgUHi5JTTHajkh0MSI6DoFfgPo0HdS5DNfl6ecX33mJbu2/V42vd11mPU1G
F84skxcd6Z4IBemxUShcgC5fnjBF9zd6dfrrnUViweiQ1ofDnDHpzyh8T69VNAw5
ziRWNV63NcQyZCMdzu7IRgbAFrCT94NfU8ekbqhCy5wR7uNoepXDpEx2ltrFWFJL
43PCn5WouG6HLhD+1menpDVDI4sn+W6KbqIct4Nf5VvJe31ZW+XUROmx8evkmroU
xSoCdpSbNJ4uJfk4znl3YCYqScJjm1y8kP20Ov26ntetD1WCeLGqHsp/RRmS+Ela
c+uB/3NshopUL5XSEWpGlH0Pj3g2W1gdGumIzbsArTlddIJlmFAM+lCNXrxHZNBG
YTGyDgeMsqnUhQGqLs2rLpTC7tqs3VUOza0LaLfr08QM9sSqCPgpvXYkdDdhTM3q
Z2Xj47xAKoKKMKt8b+OX5daDalqgPdmPp9efOdBBlOJGZFkKmUKKB9jZQtiH1vXI
jzE6hyso1nCl8cCQvKUq0vOymRa76Hn1VKUQO79yUG2qda0ml8eEuMoCEJCsvGuu
Wt63MerZCU1yDKZo+U4fdb4gOhPgkSJCou9hjHWjlkVHwi1wz0WnLk3Z5g58nuQW
Dzz779QgvLC1UWssTafVUBIHMZgOqHl119c5BkXi9NDyPEcAH3t7ade1NTGt50Qj
ZauDQMYtLETleI28qUMIomm+ErpM/I1pxVCQHnejkKpqYVIgRr4FDjDSv+mQS4F6
2j07At/bE/frMdVNdcRPTqmXWIq1Oji3toNUm7cSs5EJfYIMFMPu3N0zyVYgLfGA
vd4EfBu+Czv9bR4JlLZcR54EeAOWc63LpJ9kd4WqQB/jMwsABgiG3NwoMvrNMtgp
oB1ALFr181V1ymxC46OKJjY7xER/9CTbecp1iAp40MDCdXkBp7rzDeIp7qEFSLj1
gEFGlIYIe6cGUuerqDbfzOTWdBYsXx/z6k+dpToAhI7lgm+M3MuqySdEhgFCTEWi
FvzNaJNIiIox+NsxGt3nBZvF6ZhjgXVQsjaVXlqBt4s/M2OHDPjyXYg5dYP8Syuj
zqlK4XMp2GonW3t7H/cnfxCImHg0CiojUcq250owa5GAnlHvxnxRm5eG0WOe3X+s
nOHZoSZ/hc86VqBBkK3uR9XLUyAPyO/xadJbWcCXTmdFnIBzpgbBZn1l2HMvRLRw
UGsu4t/8BEkKRUk/rskIrDfI65n1NQ7/K4Zz4729phE8q0NDlN/lm7pAbpDiypWK
s1VGmWtpGLim4qH5eQavR6KPue7ySvOs32eT34t9j9PDq0gAqGHnB1hirxSDG+rJ
aXHDbbDchWH4bMmiU6uCWjw5slPqL/DhDQHSmp9bicqTLeyHsv9sR8GbkvoX6J7j
RibdUQYBArRM57e0Z5diICLjCtCL2QlTNJQyADHt+Jz6ecaqWS9wErHFwbUSxKGp
3XKd6tzHWdaqrxwgiPhCrQoAO15rIx5Az9xD3tSlj61NI/AdUBpBACrQ5WIiF8N4
PuISo+VF+BYi5ycH454Pn2DHu/HVMNdbVFSryo9o77ukF4LZtgkYFiY14qWkMdQ0
/Ubxcybg/ZhZROWkWReVm5SvJfjNVtae7gFs7u7sumr14ckehh3R1vJVSnZi9n2c
5N5EL1+oQxFX31nJNg1Fy+afeXurpeascx7fsy0BaErQuh9u9fYZfFXWT9lD9kj0
sFKsIJyl1+4pBOytSo6WoB995y9yUGyOg1TDA2aaCfCcZMg2E3kZA76FLhMxkBcE
BPJmyhAe0CsgusW23GNgSORmVJjMs6aLd4eD64UX2jGpyPKLciQmTAuXp43+INXr
Kp565RnrwBI8ZnJkY4YvY//kkfYCpSSJL3tEsx7w0aVYQEnY2KazaZu4q5COmuP0
Gq5ies0IG0zKO66CYnVfk/N/HFKlpm1idjW1bcUeZ7Z1mgFMTSaoejWA8zVaU3Z6
xkZ2xP+JOnGXijqWm/lr5zjaJABjs0iyUytyQtlVz0e2SEm1xc01MD+p72TiTXcu
OujLZQxqFVg6iUDGtklrUMk3VHC/0KlYUmLbayK2Cvz2GidV8yFwOKIPLObAfrtG
oCNoTHDJNK4VUU1VjQn3A28QT7sNSCWVNEfXj31D6FzHgASgsttStoVxAdKEvfON
NGlIZDDDbfUZzNxwIhYRG8xXZQ218F2/mw7Te0oFDDou29VSrFwdTLjDDKOcXzJw
G1mBnLPOe47xHjOovp9SHlZ4wfzwtCsySDeBabSJALjC9rUBYuv3SIxIREUVNgpp
2cTU8G7X+kSpRZWz3TZvSpxt21cPxUVe5n7TtkygdG8Luk/5h5amg/BirzH5e/pe
6Lkpmf973FLbgD6Z4Ws/VbPw5SWgNndjubT3PCifvz4gMzFlts8TVSfEqSVsx+Xp
TD5lPKni0zwh8SsPVOPqv9a39F9etgbXhAn/Kk90pZRQx8MBidcuSG8d3tflo5KG
bt6apnBlSmRhhP1cPwtKWx3xwcUEeyp69PLJU9ZMuGDk9kAZu9aE778e0Kx4mC3n
NT+xOOaeY09PSrthXd/dYmmP+k5zGVMqCkMDKMDL6mxicflJ+WPgxssz1NLNV75U
xkKKpo/K8++X3Do3uikn8Mqv89LEHaIw2RZVa49in1apEU/a7uwoG7HuTf2XqYTI
1d+Y1XFzrvjVDf+qjOMj8BkFdLx0nzJGXc/dlJhkiy4gLLRnvdvjPpbqg8XJu1RS
YpMLASRKoeC2wo6YGAHoTC21+Fmhu4GW2HMuUv7bx/qkETz17r0qNLyBjOFxFtfh
pX/g79hUEQYBsltbphectvCcXrCJMLMdnNjM+HbAlF+s1zBEFpAINdNagsOeVDyD
oCv1nCFCFOR+lbKMKxrZbOW0xvvlZZBX1rXauJ3YXYAvdoxqT1ENzSO0O+vLKs1U
j1Gb4Kvh65dscbJtg443Put85vP5P1UOzuRTNPzguZcn0yngsU1Zdkmyes7ZYWS9
gRgsXeEa/zJ0G87vG7SJkmgt2884zhiacVKWGGtUDf/EQZaC3SbVYQZ+A6DBDcOX
EZzHQHqKDBS49wJFJWBn018UDwrufdgj3+F5P6+nqY8yTxOL2UVWleKG2nqyGGts
12bSsNAQuVZ3oifNAFQoRKBL445w6tQRTljAwVUxmZE19nHnI+bPJ4Z87CnODq0H
FrtJmlEN80PjjyRTLkMYyZ2cFL1HzbP/ckjjKXk68jh6Qc8RNOTA3sBB0dZqUARQ
RSm8R9RGW4UR411kZTRXQokdn8Tv0jkvkwBk+JSAwXizcpJbk1RITG5Tsz5C3rR5
aL/78ZS0zmoCE7VwboxB0+1AuF5SnCS3cKr2aTbGWtsqSEWJ8OJDrX8XrtmgeF2p
pQej4VJYBttMOFaGWt0YObGDnoiJmX8BiH3zJqohgQu4+LMm4Yvl9PSib5Q4J8Te
iQHSgO0YIqdwtPSinV/xAvL9PALW2U+IkojSrfeg0T3ObTV2uGQt6Fqkv7eSvgx9
TChNiewOD8r1FCodNCZ+JU7b/AcubHuw3QDTacrewV9Jl4FCUnxBEL+mfLTbK7dt
nR1dwdv1I3/muRnCG0B/3d07gv8K5sl6PFXYhs/PzucdyseyyKZhFk7/71W0aGb9
/s8tJBqcp4KZs/C2K2EQbkqI0eKgMh0CFjdbqTFhWmb/szVplDA5eBOgiAdCf9zg
zis/g2FG3uEmm6yi/mwIKdeh33mF4zaC7cOVaSoEl/XrMv3GCzvu/J8oYzciYeBf
PXd3DzEAcNvDZa1eVToZ2w1vV4fZP/YWGREKAbhD00NiLt3crn1BgtkuOP53JAw0
EfgbTecnoQNkrPmjEH9dYdfoHQ4WT/VAwofqhQg+9kOCF7nUSg5KivGCDXNxCJCf
bnrY2jrXk7r32fY+ZP9SOTTLQwTtrFmQT6/6TJnIQoMqUDAM7iEmAZEUu4gYdJAe
tidkG5xBvJhc/SNo2iTF4SQAD2O2GpLgt8YSF18JNFGlz6W4uPX2ml691KHtWbpD
/3wxGCAEAYcmKOk4Of952NiKVGn66i5NNb6qzdrK41Q9peTDQiQCxo1CtIB2VnM6
Eg191wseXldOPQPu4ciUukpmT4eBGQqdZuoy0HSpUU1jutlJwkIqkioxnN4X/wNL
TBBMTRK6m7PyVS73jvvK/VEfLFEYEkWoNDVN3LHHEth9roQqIDeNROtADD+uiyIr
uusG80B/jXDEQ66mqzXvKLyEkI5c1rtcx+kl+5+iMgKcjd8MMFEE6fwlK5jr/Pwv
BG1p/R3r9xT070AJ1SP42HUxSY4xNua9iuL6ftOjMD/Rnr0SLIMd7nUCk0lqw8ap
1yA84zPhjbuvI5piQhc9sjmS9r9SgXAbg3f+AX0HKmuo0sIs3dBJBSMjT/3csveU
krDrtHyCNFocZbFmzDS2+m6YjTrbda/yODzm0/V7qrpmbLw5AYUniOk0cbr/l4g2
efrDfuUrSdUbzESOtEkv/Gg5e0TYV2j7yThF155ZxLTMqOHo0ITOrxsB1UDczjVv
Ff9Y9J7k8SKwBTlImEYet3pT6FHT2P4+6xMeQ2sQTZ66bpeaVxjGs172rOvGoVlH
hvq9lMpOyk2r6iuX04SkRLc7MlgyU1SQS0iWZcG04atrUXH8f48JOzuU49gEJtq+
mnayaMt2J24XjNBPrkWmdOB/QM6FIL0sMRDPklqsS3TydnnqRtNPVtJR97lE53Ie
QLNC9sXqcSaClNymwS2ERdIWe0s/6LspuMZTw0PZ/lkIDxSSRx42Wp/HNn3IjP73
2AtgCh7T6eca+dt+Rtx//aVE2RibkeumKWj9XMAbfDK8FKlBlz72c/xQtB2qSzhR
7QsmSxOxzYRghqSFZSA7Vz+oJhB/pB9/xdhCIfUtgxEd8xNwjOV8RO8gbj4j+9Tm
9g5I6vjTYibI4xFU8w8d6ZnuUzw6XnoyizRyeuBR24kC5EbJlydt4nnPnMIsay+t
RusqlUX7ZN9DquVL8WJ/Aj5O7lOAxZTo3nEV66UmkjREb83aQAeryKaVJ3FB6U2e
7bEQucPPPvEN4D2o9sffNP+kgm347d7iWbf1d/Ub/XjVQ8jnc8tt5P9RAnBwUtY1
EYIOGqOepAm6rQHfhEHUu25ZnsgbNQ58cLZzDcTK52HetJ7DDqVCJ/lZt5fSTO8r
BTeQYFy9vMI7jHQEby9Q4ImD09t3y9PAvW/54S6PfpkchZ4X8Zwm3eq9YGtgpyX9
a2eECXUz3YiDcevwloFtjWMYE9NMn7K9+b3k6TojMAX1BDFLw1gaE7P7rPvCR7tO
Qwi3OJ1sTtoI0p7FU/o0rU3oiwgXbuPRdAzDETFSypDoc+aLsjUwFtLj8N/8Pvtl
GZ32ZgPS2fjKssGPSZrP5jlB5SERGQ8S8fQLuivZtzLFMynncf2eTVKyviZe2uEx
ZH6V1steJWbTsricCAQ3Vf6Tb2usfS2PNt6o1NKtMPvwnTOXa+rp6dezDWqGT0Ja
y3o0mEZK4tEE8xr+V1jaoTPBJO+89zC+XijHPznMc5dg2KIufo3Q3XROFTTa2W3U
1wsNeY2bYrLg+yqSs3ihTQee0ciMhADBlhK8QCFzdeWzWsoDzWKGomzs63vmCvQG
FlzY1xyoSdIab/a1WQrjgtaXnTqZV6VryaUpGjsvdIFTlV/we5ukptubHtESAs+i
L5lEAgA+In6l8uyXlqVSo59yFdOVZ+NlC/Mv58soylr4BGskDhULOnE5z2qQKtym
ZVt9P3v5MviQAeIpTbbaRyLjUdDY6OdJt76G7L8kqAycuJISEb5t1FQAZUtAx9xq
tehtsWh3+HgPVHhV7kTE77G2QuHX6lm2/GY3183i1L5eIRB6MAgP2p7k18oSeB4J
Z3dk/VnaYk7x89KOJ/oUmcnT4i+mXnpNSNwqLSHdi9ye3mpS+sMLn9ZbPpaYNlJt
3Wbn4j7kBW1on8bUEYCr/BqlMEF7thFB2CGX7dzVy25HXXJMU+AAzFigaCRlqSzW
1hMYyq6GTP60bIwDdTXkalIXqoFlFNAP8qdmyiD8raWqZMKPfYN5O4tLqj5a0ENA
mU/L6piehgu65+ZKSg4uS5Qd8cZgLsTXrcP8Naa6TRQIUA8rKjtya0FfUJNCZz25
vrofyI17Ki7dBOoLCJRHLPTisWTaf81fI3uYeEzv5V+lna6ifDT0eP/jXNPhTNGi
jiJ+Bq1yieYSJknxcFL2awTxcNtUFnJnZO7tqFrt0ry2W9R+SVdbviPXzhipHdoi
tZacNF+jKDIh38l057hzPn0z1MdwQqshanFIrMPTx1NKFzOM18veLAMxWBE9/GF7
6CvokrDtD2VWyuTTiOywL02WTu6Ik0VyXZA/8f4N1J4MfeweQ6Ggjow49cpiU9MK
xvJbBIOtvWyjsnvtLxnf1YciyGplJjdwTwYa5PeuuiiGU0CcFdnR3jgxnRV7QPI4
ksaHQJcPA8u3kQHWIKhhcFnHCNH4uVLkZPRxq61Zuz0rr3pEFjUlLogxrPH19nYT
X8j0yog+UQ9o2kIqef/t2JfATyZU74CzbQ5EjGtCNCCUdaHGJi+8Tygw1Xvc65hw
K7oSTvG6HRA5bPn79jGKtybztt0wfPpoT2Kj6NKCJbNN1X8732MjmB0uepl6sWbS
CiMGPGOY1ZjuyNksKQFGRnosd11y2dadvkR69BqK1izVcq0lilEU+9CrhwAJsifb
vIIK+C1o+wbXUDfTNAL/REhJj+9d02ZGV2DaELrgHX3PCUDzv49hZWmrI71j6KCn
T2xfBfljbrSgaqMaF9CCKyHh8xTDtCEibbAiDgKQmJ/GkbE72nXtDRoQebm4ZS6p
wSsMmcOrKOfBJclcv4O8nwT20t37fIYl3DFPLb6R17YfAbdDjx2j7PVznsHySBrU
bletosLPDOpja73gcAYNXePXRExrj0nAnyG1mgJoY+XeUW5wf5rBkxw9EZFdzxUi
+QZcqOa/ThDYIXpBAMmxS49Suq6AZaGD2EgJn9cb1s8kjZV13ydZ/aUJWC1Y44wx
mcz3sV2DLoSFvA0xEyxbmn2sHOTrA1pGRWJ07xEiwX1Y65/xtZVgjNEbxdlRX0Gc
vDq7wL6xVTsI1q1UZxVR6AGemZzUYZMqRh0XlfN9aqUnSUtHwUKs6ln+ShoBjmMS
fDSPsqbvqtg07pAr7iAcuMg7e6c7EAbTfo7fB+QnXCDuLC4g/8fWPoFImKI7bSfd
xdP2A5mdxD8U00HlseW9kFrYBoVvGQxWtXNJvW2crL4+udbcfrj/514jv/mONKvG
EGCxMNTqoCYTalI1oMniE7foBGN0+xNPvpfMsoy109tWvxtSbmuvuKM9KL8sn/vl
qM5YcflnZmNHWoc54gzO0wi9qRQwshDyX56TsfnZRl/lZMP4Sj0Ygtd1D6iRWdPE
Y02Q5NWM9lK45RCAu6YgmtUKftdKJlbxu9cFEBzQxnUI/6+lFpehApcTsifbln2w
tFTJ1kLNEnNe9ywR8MUuQDib4rpiuxsf5uCp2+fzRRDDi39N1kpWqwpigeQ0Q3UO
aIQ1L2WJNw+O/GwPPiV64D6/xP+qDQYvYqtUOpNBD0JJ+1eTUC2NScUvkeztuXNW
6b+4n7BqwVTJM8yIMGQbEVK29vSJWjkCkpCH2LByLLOUpOtU4dW9K5JG23FrYleh
aSfp7g4s3QL4vhns2yiuVlfvFJQEssCzCGEaElUPs0eaY8qGSM6P83zSxdhiwyRg
3RCH42sqCaXkyFQOetGjlxpG0mvOpVWym+NmDmREy7y5IMK5viRlnjX1rDCPczQ0
DOUzpyPtbOOBmb5dY+6YbpcWLWyp0c6WnUNfTlatRv7MPzL1gWqFcsf1HTpL8JOs
EfUQDSgeOLzA6hPER2I15//7vp3M6t08XHysMSHKDN7ITceSFM3zhxe9115w+d+T
l2GxVV+iPZQbBmxNFuEHLvM0iee/+JTsZpDAQi+h5MB4jbC1hbl09AZuJKf5zpaw
QzE6Ev9ngoYgsx4PPiQIenwEx8Stpd5hkUZFDt8MIgLe1YbXOzv+eMdixr5YvkXs
MGpsHJHf08Nhce9gLFACC0pQ7epdVBfCMCnm+q+ZUfw6Yg8BVdBwkWP5yg8/GtH6
ZVbPDRO1fp4yfC3gMOhjjGWIA2PKUy9YJsNSM6fCc/umC55DNdyv+g2q/ceREV/j
iO72inrsvkOIVf+tQOO9R/PbPB/fcN1/nqAMM5KZW2iBCluR3K2N2yzPWG3aVIJq
EhqHIbbnLjVfn6fy54lhlNsYVjbCvIGBifTrw4+rk3nrH2OYOydenVFSZDy5TmYG
91aNb0aR6orEyKPqtQKoF+2HdffcdhkzLTP0Hqxej6Or+DtRffa446ZChRTBtshD
2YN3BvsLXM2htosh7AjwSvHMu6dZoxjKC0yuKRzQlac6DlQ4F7M6NZ+LUqyO7ycA
H0uf2IttaKFH1HAmG/9oBcvtvPbIJzg8OUUzmOoWVrAY383u72NSQH4uKshxrmzH
r1HpaluAxXaf51Iu/T7Rfv7NJwlpnk+2/o8pVq36UYGFLfMfdiiK5gmRPwIuhQVF
CrX7Osq7xRv+cmeJhkXkWla2tVSeTe6ZyHe40L5uXXFTF+a3viDrpnjRw2iniiiz
iyU+3m+gmBESVCgTctaB4xWcCN20zubLp4QUx0WT0kIjXo5YGZdxcNPyUlHByWA2
1AuBwnDANdoIMzb4sM/U+6a1GfRvhs0TPQKtC/n4xvYw/0f/VDKOEiIJ2UDieLz8
Lfz5uPdr4AF6BS3r20ESdWs1aE6rfb/T0pWRR5RNKVEG0iKMmfdQMV6i5bvUrSyl
h6Tp5LUMaFxTtrFv/wfz1NjKFL+0zZe7RPCt25ySKtiPQr628/MHK7QD6b+NmhXP
RTs5SBpL85FKPTKtm+Ybzbuc8uaD+wj+G1t+qj/8Xoa5AL5WpWiDSfOsbx1gQbDx
LOREjdWV/L5vR7MO5Lqxe69m6J8z35Lk+6l914Y3nNO6YrTCbiBPKPLS4UXb3PnE
3IF8teKFUCRQYIpFhNp95GYfSmJ1nNKPyHdlFPSNzf87QnJzNxvRGACuFX7jPDKC
EDweDGZCmk6iU1ngKL/71zGtHhUVyymPCkAkfFusOX0Ts3D1jYr1sEs7MlJEb9WM
/HMih+PIDwnqdolkVFgfk/egJHKGpU5a/pSNdbZrqINzQchCAGd21dqAbk2VI5X/
Pb2t50eHjJhu2NChROMkuVmbZSlwZ1I+sFcHmdpFs2vnbS4xh2BKOdsn+KiNE7tg
v0ESAr02HLHbmuAGN/t5RozViFzivJfZZ3ih5EeEWG40XwcRKW1jSmrqTdQNgACX
fhSOl1YppoE+vxxIPJlclv7dZEsSiXiNdMj2k2odWKrEpM43zbNMsRpOboZ/C+zT
n8E0GJd7wt8IPuxiUVABFXn41PdU7N7v7NuAkWKArEc2m9rGKLc0581mpGOdIh6D
HefcABxG++I6ancvtOystffFrvHdSbs9LD0V5IJx3/IDBsvLJiu1+NtYsF8beMFP
O7rwHyrvE/j2wInX4bt8HDe+3YkM2ahJa8Km8N8QgUfxooDI6ISpovdIRoF7q9Bo
CEXvNTp3ICTL58jUi9hGev+JpgYO/Go/1nYWM6FjhnDq3pgYRUJI2fOtXOpcyBxU
Z1ZbqM2xPF74lbHvTneHYnoDA65gmTgUW1X39IvtYqoJJoMELoJs8TFn+gyAWsQD
u3KAXPpznzAYLktMV3B6lLMm62VGwrOk0oJu87G7h5aSf68cx9RK9ZvrrGH9lqzA
+aD33oBb8tQlIIzSGAWN9iQlIB0ghppuJ7dn2PyMX5kXF1Q+BItOJzrk8bq4GKVj
fz4ekGkORjp1lcxhgZ43o1h5nIJVYVsiqpxL3xiOF2VxPVyyHtS1Iwr+J7Ka6cSg
88o5Ld+YWdBSPwmV7PgLv3IuPGdrBVgu/CxoAmZ9QEOFAc7iXSWXZby9eFhwHV1P
1A6bdSmII1+e1hdKrLKTD10bvfzSKjCvbqmWi22QtboqqJeTeIjMydKJAgAvMOnw
z4aR2pBpf3RQwDtWE3P2oazDbVBjvmmoul+3vLGUwZmUE2MDWUEXCpUrSHjMwqcA
uDHFQ0Q5wJvB3qo9mB+13tlBWdEZdbtvx9lLO+a36TVuLeVWISTnZRC5xIiDxih2
Nhd3yg5xQgeLYT+6d5XRK1INY0KrI4xKvEUJsCaGolbY95RxY9dhE6tZN4g2b/Tu
qMch6vMU78MCkZvt+f7NDX4HRukRoAFQvh1jk/5mGPGx9ee1KVZ8zbG845lbAzlz
o/AEivYMXnWLtLQHS4VYs6LD3BmozKK4ZU9LX6YJKE+qs38k6bqy9vGxR/yGNPnW
LOsZJKZjs4it0VYCtwjVrWjGxI5cYmS6mG4M37BuWioaNLu2DrJJisMdz4AYjEHe
pxtRmCFr2t2kXdnUKlIEVFdQgdHvu+g3SercFChft858nLbwoTISPiWGMCyBDFW7
fPQlcWvmxBYtqx/LLYQXH4Ix+Z/nkX5LS80MUOVEOSjb8fpMstug3P1waGDDosNV
pqy2awTfITz4ZS0SmORHCjBZAzeXO04Ikb2S/F5ORTk68cNC8/BSfvwdzhibXi8H
xRrpfEUL1SZxgUO6tGMUdotnltSJPlVt6fUUW6uPBWQaFSpxfYMNtLEayAadi+kv
oOlNVyZiYWHn/ILLB32GNm2ijgaKyaQbdVbnklKPrps+/V2IBBkGxHy4cCBzVUyT
jDp46vdF9nEsnUA+LUnjowF+ZoCc4NmeXTZE3w/eduktQXqRCNOI63nC2ZP5zJ0f
mCRnL1xuektTdPYV296hG7heI0RXy4yOGPes53fYP7JpMhJ1LYPTUO2MxNuZe0Ye
bbsbcMTdO81yqJvUytl72YOKkJx9om9SLt1lDl7Hlj/O8eStmlPgYSf6AZiVoLuH
/MFqUWmStcEqGwwDZJXChTvJKmSzp41hWLHwhxhnDPXLpxNOmB6lNIsCtPjyvXzN
4UrqXDMxaADvRxP/jakc9gYTt37Ingmj69X1S1mEMUnTBcMiqoWlC8eFWHF5p4aG
zs1pagsYMN/mC44i9U+MQqnhL53iya6zOrZQ0tSmC2uPqUWosxZXSIOspHhclCvi
yATnBxwTouwZC29Eq+Fp3oT4tsKlm1TRH1inqzqCxkueSZXVowzaaz3olzmfSFcH
Q1PMSD1eon/bFvTShf+GRR2esWAhs/yp/QAgI4xayUe/DK3GY1AJx8/v6s75wCSx
3omclWCUt3Rv02yyrhQxIubg4UOgg6yjOU/ulVtKATidHcRFMA1T5WsIvDT2gzmY
sGGPxPfs95ykOUdoG1ERKic481e1sUTjr6Y0h1dcK9nwUUxP0Y3La4mkSUfdJ8KK
rHmbJz7ddYsBwoiDf95vPZUjH42SVO0L4HNf6D50WM/m5L2W7PS2bA8F39oHy9De
oL9HFlZ6enbW0bWCbN8ZKHVoTIVPg/6gU/4b1Fr+7myV6tBTnxrvPuqD+2U3DUbC
X3Tvpk0iBXXPom4kTZ1S/PM6NlJN022MyM0FzafSqzM400aUjN5wg5z3UbflpAV8
6XY6rOAKj5Y4masYQzkZV+qbbSqwJgyaP1dyDydUoYWgRj0AAVn/noKgvKs4Xn1P
HuSGBJOGkcMfy0KRKxJR2aDw+9xA1tQh3pUohCJLVi9iF+Chz/O1n1/oxnsEtyO1
KVr+jKzMccW8Tt6QOqy82mOLs36Yf9bbN8vP6zZNpfxeciZSUgi/RxfYJ7HjTIqK
MN/16wW+4kN/aqgE7WRWuplhBTtiPWYDx11T35dzi/Q03gA38U9YWtBNyTEalhk5
h117p1HjKaWEsvjNAZpXVKbq3WmeQPsuJcwJJTAMcW+krp34TsOLyN5pzODAZON6
CAPCXMsfg1SS1OZWrae9GznZaUI1hKTCoLr/A0eEhv9GyfV3WoQL1aZERjA9/4hZ
t9OuU2wl7oJkSwNU+Tou22jWK3NbL967d99moz9NsNCjfKet2XreWfY7+3xX3EHS
e3bAWz1ypyZfKQUh/B8Xmtmb5PcMHkyoB/Nl3OCPbSG8wGuVTnk70F/5t5HPBQlS
FA5eZW/LpooZYQm5tHBd7UanpRBKrMGi1QIB+oO2YYz4ha9oVZy3xANRQXIxZbi7
ONr9V884q4HgtvREEpNZLpDOKbqhn6PyLHQxLhqQt+mCUs1p4eQni/cKLehK8g74
7cwXFbAxYL4oZbzy4+7BLGguSYl9i8sVR0xZEzQHlQ1uLzcCTnTpAQckg09ZI3o/
+L0w3Zs7sHYTmUclwrTvE2fT4V8WTat3fhIlDBVTwMmgZ5jaL7e7MvJEeH9EpZqE
YAjzbSd+iOulngi5fxm753VHlN5IGFMJ5Al0DGJXgabctJwkY9fcyjxT/MjFI6Qf
5sba7xKmJJ9MUfpY9Zc4vC2QE1Cdx9eWq+6sFmsgOXIm2gnEdboxrGEwHtKpT/bG
/qtibCdfausoY8q9zzdi2Q4CRgsh7VMy+iXiJQlDlNX5iT1kq+0J2iEldehyJK7l
Sc7egtxlNb9t7fBsDUB34nWJ9/mAogucG1kjVpqjBZ7YbiX7rwu3kbZ59xEDJXuT
U202clP78rjgIzXgEeoPyJpt/7oy5Yk7MdFB7Q4Ekt2TDu5+feQl236gK6ajgSGU
B8yIvZyJxnzJNYfEPBpqZrTzZgOjBk4U3s8OlBi6v1b7dGh72UtOII+wxkBDpriy
wys5o8mvGUr5bbQccdZF4OrM+ParTi2+gErJNoHj6IRAOhnvBW2rO9H60GWMRVK7
57ujNxz5zhvSPjSl5NkPCBcD+AzAZNDjE8lOQa4P+dgG0Ey04a2oPfmX8vR3wSvo
vTFDrvl0ydaqc71LOQsvbIQ28UYzOQnyh75pxGKpBRIliN0xBzZd99aZDo/dQsv3
DX15/Z60c+6veXrcj5ZXYGFmIdP90OjgtoBoJslHnKGnETO29vnHX2yQSUDrsWva
FaLXJ+YUtrxav16spX+dCzxhWyAKUetPnU9+KywacCU/GengJ1W5oSOAp4AkU/Ye
TCaBMMjmaKUFEoJtjpG03HASrrVZIkenvhyXNSsqus/+FHVy1Sdt3eQyGio+CBzU
dCfne6PxGpE8cHSXxBqUAhf1rz7deq0/nljJGieCped+WInUEaDcEC2dLgpan+DF
6XFJgdf9qBwEfsU3JBMg2YNjeJc35IxAR1O6P24CrMwAGqDzRcjjK3i0KkZciBxH
QNVbVYAcyljQZFDANbqx50GOWnv7Cj4sW1Bi39ODs+aHvBjzD7jCfAud1opX+4Rh
0PUijsXtLeLWDHk9pfr1+qWm6jHJy9KoL/dD+C5sAOftiR7bamfXvNJOkWecjWRF
JUodu8fsngtcg82cawwSNycnSZYIE0cKONye6tKX08HTgL8CzyL2Vf0gBe39BZiX
0SJ8kpGdIwveEIDnDWAcfDnWEpUze4ILEXEhreEk1GTRJRwNd4ccGF9L1+vW4vnR
1OUjGvIhfpCaKxnbHQPHCICy/POkBO4XcoOhmRpPk4JgLN7FbJlnkbCzEdMmHrkb
ZaVS94KcFh361dCp2QdjAYX7BHQWoTYG3stBAnizFfvFsrQr6TBg7LeiruNmwBtO
EYYualjkj2dsEi62zDN9HZyR5BArl27KjBEEKqWWJbN2T591QTwn112C9nUvEtTT
i4jOMERptrswkA4Ck7/hTjDm+/wW2B/fcm8VhzTcR0qxu83ELgKN5HE2sAX8LCEp
dLTUM0qgUGRFAUZqeMD+kAIWzilWF8bm/lXKSuAuSioTuklBtRJ/AzbdH2sI3ZpL
xdZqjD5BC9uUY9SxNZDitpcywXmwynCN7xtqUEGHnfeP9mgZJcn/a8G5fI+bEmAl
uHOCawHULKRnrZOteTQX5oAW+St0cikzDOW7RCYSlTrfEIiEXRvRj5XaU5til2Ei
jIkMf6OT4fuqtf3ENA3UoT1UUUl/lU0Oi6FkHI1xQQ5Hh0EEWm1Vt01bq+8EUJxo
NAiRbR2vh8leG1y5+9agBvUTTtqtalUayA5GfCoRK1kDPk8ViwIwQTAwWVAL76Pq
wPOButd8XecjS6b3XDDDYJITVw0+a6Vi7IhE6ivuH/DOg6bNApa9Gs2hTW2M2sWe
a98yQ2dfrr/EJW0WJSGE9K5hCI0ro3Mqy6OZ36D1kYPq2VG1WRPvgCQnclsQCU2E
hsiWr95vKlzQYJXgUp7pfMynh2PnZsUNvptY5eokTtfN7feJcnIHOgnclIO8QYki
AxWSwJa5YvJJ6zQYm20Uh7gkRdJVQQVqQ5OYHLQQe5F6MJrUChVq5ml6jPx2a9Bi
Wkmal/vU3/nrV0FLj3lzGLAlvVV0xN1bb61gThn7dHsM4KqUtL84iyzNhOPPXVAy
BE5yahoLiT9KneQ1hGTyKewF0legWdWUnQ5Yf2BU90iPz3d2ijkgKjG2zHMHcjhG
vMyt3AZLrtpZLNw/Y+qw6vSZMHHHoW5j6o8H9Sh48ueBeXUcL7aZiOollCiU+jjm
LF2LH4eX3yWPmzdFJhI1mWjGiatH+XPlGll5MP/JwqraGHrpe2oDbs62WpbObE2E
+la1lESO/jGBfTlolmUFf1QyWx0sDaLgu7luRl/FCwc07Kj6r8+jyc2heUiBki8Z
XaNNq/q//MAM6KiSHk/HzxYYTFVNyyQGptsfxawnhbfzjZJTpj8AyOQtqdxe824B
8Dzq1G5NnctgJHt0MBvUC6z8GJwpoznwjurerJe0peykDBuTrAAmMq2SkjyHZpik
nxxAM9Fi5rFji//yhDgG3fLR4JLqLfUiMhhnrqhDazKhIm7YJINRpnh2EL5YYlt0
Rqn1mZqg1Edyj7+735JljWtez1J4IwJWa025m5ns9Crue6yZ8cqOEqTa02MdrOnX
4wEyR8n2YHIjsOadOgA0wcZt+zlRvT2Yw7Bnw+Jg+PSGGFwCcBI6lOkonqgaTTlH
hYAARuF5yW/a0a4HidiLZTB8ZLnGKV5F/gJYHqk9RGJXRGkd1vOWGAXEIehWJKX0
ywQFHMm1cxY8UQCC1jpuIGTXK3fYs7OfxR0ZbKGWDRxRnFQSxEtkuKvnvYyeDxb7
xUjO7Bq/RXuqddgo1GCnzuuADim3Tb55ppiBXvAbL611BdP4/4qLnFn5OzHUcwxq
4xXSbVeYw+ikKL3MHJ34HbSiFjElGenSbajBInRU7sPmKRPKc6qw1bHIdMtpkdvK
SPpjq/0fx6WJhStTCtDPBAVVMz0t+n8hewoLvMrH5kWFa4iCa0gQ9zg9f9Q27nyg
RsrR7VVT745YcKpl6CNL3Zfq7bWEQNw0LViwnRSp54rhH1Kw3zbxTsGiAsdEppmB
6cyKIE69QFgZRayICVXjoNfv72Bo2SxsMRjIMtU760PcbtMbaceMwlmqlqJR92oD
J2EzRmfQMCx3EWWoB/r8sMGMVGRz3LZc5SmEDEtWlR8dejT/MBP1mOj3WNGqGLE5
oFkVFtxU+tZTrjhkUEhnuxBhzPHCBWNVqTOHrXEFAnZPw9wnDtuIXiqlzq/ZpwjX
s48EJtl45hKKri9ioPHRf2Tq/efd1s4S/4MbZAjD7VwUwBnNKXnagAM2APhp7Cml
+jYmfa2gmdjWwrqp0V9YCDMQ2TYIvkmXY3AnQvVV5PRYiakKLRfqCbJEE/qwg+Vp
Vv8Ya6kE/eLaS/++XO0ar9jukMUP8LKF3QG7ilfYTtuzEawU80b7fOPXlMv3iaaz
aqqugwMKcIIB/KxTOLv2zX1iTFqwcfg3cCW1/obwLj1+HEShQxvTF+z1KjDktRa2
6ZLtdooULF4tzz/ngLo6va0db8NeXhRONPFfRaVH31nV+a6NWjVcdoXKyfh27PCn
d6gts12lY0Hin+ObQHsvFY1mMgBnflR3wS3SsvqALYoKJ4A0DhueXXJw6sGWylQ/
YPhJCHBA+ZGIS1VoHWAaMNrl1MfD+LUzJ/95b+aG9icI4ulTzqYQOJBkHxUtFJI6
icCX3PeIQCZ1Lf/AxNHQxCvNzRVOMq8Fk8NkFG37OqzefC57HNAbmneLzu3XGAge
4p2GE07kCJ5ZruqnvE6vcvl3wcn6KfBK8/TSsiJBfQCFtxuPVDrj1J+slVhtYeE1
6cuktzyXOiiB2M/1pJwcyO2NHghsWBUiLBHU9ceQ5u4pa6kDJ79Fpef0Kwm4A3sI
N3gOTrPsJNAOhT6Bw/JYxtFQLFxfPbwigx9cjDWxepaexCSE4+KxhzmTNUh6lFvd
7qdP45vAQsfNc7oaG7ajc/4NsFcU6CP6Pqc2s+BI+Onim2yxpCSZzAnTVG+oQgge
Sa2QQXfwtQuiKJYNnobwfLTofhJwFp9Kp9T65ZLdqLNiUwcpxs3bqdKAXD/kx6ie
WqjjtmraoeJopU5IxH++2tShwQaGPxzjRqd8ckgLcKkLySGdzmoNBAcWqTpHAKH/
X89Soxf4evmltzuiF8xQ2y/RLSufJ1UFqQ+Mxy/2x5egeKcxPvIO+du8ZV6rW9ax
axfjMz26tfmR+VYNi2YFr71AYlTTEf+YgBMuIb61vf8QQMMhwGxD3fHWwwTSO8KV
NSeYgsLeCEbRLnK0jpkQWIV9HUPrlIRVBrcz+Mqa/D4/6TIRjV64kAR8sWxHtj2s
5o6ZX2f1kcYlqivYoIQoUSX8lxLjxmFWLUDw9uaI8bvlXfn2I/7Dm37DIK9L3XxI
g4WISaTWLbipkBxVgt2WqSU/Q6TmucnCfD9byCJuG3CMjo/RnQbjQm9JL33q58Un
ceLO1BYI1nUV6p+DPxgL+/rYIcTWvPeNgtac0ZovBqj78wO4+QJO2yTd+G7wOMOa
p1Z/THoqKmCg+mCgh5h7I7JBquR6n1z9cwiU/Ly0KPAtzEfpNTWTSR/XAh6Te/HV
26Is/jhpu9IFh7llXF7Q91x99/bxyV3MH9faqMPByuIun+p4xMspKZ7HhCTmWTHq
cM8AFKT9O+xWug9bLLp+x2vbLhxhMTAyRscGrS92rDBHQ3PfzI0NPidm5/APE+Aw
1ynOcjFkg/JYHWF+Pi65wW4uWTZNogPiUt+Kmd0pUk3/yYPsXHk/eQpnZrlbluPt
CQkQcJOz94U7ulKDreyywjopvqs8MPznyjMsirAvnwBc8IFQbxBGAvPrp9RvOlMY
oZBVDQ6TmFv+s872OO/3/o1uC9SnRVg4UNQih8W6kSXtUq461jyTTAyioe7tN0+b
K4+oJlQOw06gupRPnF6RwHvgYI/aG8p7dqsuiMM04By3lbs/jWsc18B+9kR7DVI4
bUniQpdzN+hC8CSZFmxab2JbGrRYUrQzvjFH6xgDQxLO23SymjdIwnfHPnFrPH/0
PTBQ8WXUeNUjCbN0N/IHpHFjc0RGXJfHMzIw9k5VnR/DhtXuPvrYnPS7HUjHGVUN
3Ql7cJ1KiINH8zQCCcpN2+I+y0NzohYZPfpyCZt8eJeLIQNiwe6bcEBV5AFSRQUA
kYC16WksckPaGedqkSVzoqFQwcoXO0ggf/xIIpkut2OgfwnWTZUzgH3AtFNdCD0w
LxLp1zH0bfoV+kLy/MZ5iDRNN5Wjiakt3zHvQv9ZWCjXEZZHPG1WtfcHdr8oJqaq
APpe26anu8Dv0pYMFbTxOM8/cfqqP78clzIgWjbjIYISkm70Ensekj8PKYE1aEQ9
XdtIySWAXFE/UI7gOAUNS3X1RJzSNC6iYy9J06aUDHC0EDzR0KCXd4iUkMj99uRH
v+zYWfiUn51y4GvZintkrHulTyxctYaOEHNEP/8s4ULmzWXC/1Sj36cSEJH8D5WC
9CMseIrkiXqD0NA0pyi9QZOgnA/g7V603vUPCDswwr4bMxnIadolSQ8JwiZm99nX
9FdE0w4HUm1J1Vtk42hwBQoph2OtRx2LbiJGG6yZce7R2N1FmmZzlEO1T/Wm6pr2
Y4DQ4y2w8RUGo5J+JfU3x4tnI3H+eX/SQmlQ36Ohm2NCtHhk6PuJhoT/I41YsTXB
3pWsjt7PZPNHKUFKZV4lNJs7j9Ge2St9X68CgoAV05AxwqhyOje6rusctwpOh5Z3
Ff8wE2VvWvUUzTSo0Am9wy9pA46jEhy+Js5Z6mZA8XHTIcsUDFbJhYEydesLm3l/
FuSDALMQKu2yWMWJ1z8YOfjHYiMIfB8RnfP/rgbR25ym8p8IA/50PoMnfHWDGMey
u48ad35Z+H7EN74XGXxsw0DgrFxdN3JP2i+vb8jfn24duKaJuW6KScAYgwTmiBcy
b1Fi0abGuFfMzghDafcsGlp8eKyKG8iwb4cA4sfRxc+2BtdTgVKbcwoeoXH6errw
fLjYgW7zVH3vbm0NdAm2b/6Sq5F640SEHV9J8xoYfkJGhHH+QcU8vVcN2yBYeJT6
wlA/wl20zl4SFRfcA+xWw671ebhJHpeyjnu9Pc7Il7Y/SnE4XIdBkRNkasIv0e+B
9zK/rVVc4hlFuIiy5hsJecMFLUnS10/d4YxSAkc2y8O8qfB7+SPZ45TpGOZayqNZ
NR1FTaw2VhVKW5zpYb0LbsrbmKMIG/y/MCAwCt3OauuZQRNegYQhYxkobW/KCSG1
neKrIyGkpg6E4ATnZEISnH175is14LhVw7CQ/oZhbv5zgDOmwTPoYgTIv7EhdSrs
vQ8ZcNKLIIflMk2EZfjFSf32F+qM4KNrHXtqa6zQiYbSwOGLLlMPM6WFTEvMT+p9
yT7429GaS6Df8L+eblclwpUCiuXojpBz7wH1xlvYgGU/ajn9+XIyHU4+uaefR+Kl
nwPyo+iA2gfCmZlvG6PH/AEFVOwDjw0OLTADDiQtmgBp78GTAks7L5ynEFjI91XZ
7WjGnvdzxZj5TbSbFfqTeDFkjcNBHlS7XThY2U62+vaHpt4jQWgmlVt9+xx7LSPE
xaDKOj9JBdtMPoNf+6Jj0PAqhPe6a59mc+81k4O15eJ4turzXWTtalDhzL+zyNpL
zGQadzoHQ2kIKt/Y+1jPb3hEdZKTefxePPnIItXu/0CkmCxyKwyubEDrT3zV82aS
/hIpHW4yX6/LyPZZgIhVuLwK5jYRj3pevbb0upG9hmQEFiqTHOKzCeqGWXh+o4dN
QR1T8fq3HUZPMfHYFCwl40QqJWQn3CIcaFZ1BezH9t2BgSI6FcnfY/De7CMzYnn+
gjjftUs1JOoJwl1y6jgAo7xjU96Sowtd65gt+XQQ0w3jIzcACsRgJ/sjJYQW2oMG
NkkC9q6jCkVrh/CkXoqFSkjkkS9W/QSObM26lQ42g73EURXKBr+bFLzbMnj9Hqc9
0xxa916v3B0VfAsmJW2psc+XdBFwxHoFEUTqzMBuoLzsc/DNisDOD8Gy26N3grBL
191W7B0aL4uVxXS+bFcGxl/noKcOJr+nCqwWKYyPjhzgxrj4Zaxpwh+t5ZMhgm8s
rgBEvHkMONcii7/PExfOZqV6kyO/kic0aBmLoGMleqXk0w1GWd/mFyd3AzuhCysg
4tEjl8bX/PgyjkKTEWAgxSqpPSYDq6+R4i8iUemTBnmyQNltN2XVTMpi3wdZdhBq
LZhknC/UXG0bSj190baF/0GFyHYP+rV05HiH29qiwo8EoW9qJjqBom4lL9Oufpjj
X7hEkxcPn52+3w5ikcKkvFeVZvmiLhYlTpdcy5/3CkrYcFy0iL/8XVBcX+deeuOH
gupeHZISDgb/kASF7o8fryRz/SaGenn7vSwHGc6aEgqWdBa0UCnSFG3B0ydVYHI7
MvY8dPbpx18hecaZPmXvL1yzN9SJA4Q8IH2a5CiebLEWmvZf2ol+IgRSCOCfYkVZ
+IdQLw8jCXf2PUxkYOfoHe80uV/Mg9cn+hCwr3tHfKaN9AY+DEvFcEtiTxGUXb7P
KcyhlKfbvR+jxE1KYJZbuw3Mi9aYj00QXDb/lXSi5kHFPA6sRzeHVwO5Qps5GWv0
MXxlUPJO4CLe/fDjmxJBE9Bgi4eAOxH11+xYbVIYDzDw4lxtAo9Ojt/GVeWRiFAL
OHf2/oRK9Xa4Pw4R09IHildFYaqw6eCsafKvLKH5owGFBFIRV6ZPuF3tvo1RQxX/
MBNoOSK9B7DOdaxnpeghBtI8k0mQDYOUEtIBvF6o91lnNcHJNqUCivBDOFqBKBX8
kCRPj6Wxzev1BLLLKUyVmmV9Ykask9xOLOytOBlJbcnvG9pWH7/VS3sNLWVulguK
+YpvbgCDik716p1OUh6rq09O20wPbQxrRc8nC1bPkeybfrA/wcgpAHiYGNp6QR9Z
Ph81ix4K9oOPbr/hWS6i4U45cYih2YsaVbwPB9nTPw/78Y3UdWhUw9S1X9GQmki+
+FcPRWe+Pzwz/H6rLmkYhepQUkLgpg0AvrdzZ4trvt7Q0kq2uRfiO3Gb6hnXmbJ8
3s8nY67Tou/+tcrTLxLKXbQjuoqzkCYPQEC7Tim6smHUm4DUcXYCab3yJUWqpB/F
SZ0wWQYTiB0u5sNRzVSOMad759r6k3ruwB/myI8xZTWCZfnXPdTzQaXsIckk3agS
7slH5RQ7MnYviN9x3Ex6LT1oF+NcR3pMSfgJ4py95N3KF7iEYkQUbHMh2RTriL7f
EBZ8OosJuxf8ogiTSzp8pFnu/w9cMgoQA8rie+zJUGSDohytDcgRzGIHhSXPZbON
/1uWLV+K2u0AkzSUkDSdilYMOdqKpbop1CJ4nODKZ9c4njhaQLjGsV9bPSNUeaWT
j02Vixyksj/wUflRfqYFehzg+tcherRDRsmnC0n7vb8zm/Y2OZ04psTczh3AkDIE
7Przbirjnmp/HK4c3WnDHW9DjsZOPjnq2obBJTunSzFy//zAuBeGS2Csum2q62bG
Am1dW7q1vsB8o5XqbHXE6m8oqWLKBFntzXOqZmQDYlNblP6cWEwnK4IWdaKdiEre
+bN1OWp+AH23VdvhAumelF8zfMzRp+Tm8GV3n4GTRmIrA5J5zfdxMzcuSqu75OZO
rJepNCveObnIkRytR5H2lxbaOvbNCr9ykA5j4d7lS9LPeIBwQiITlDDGwpqS8mdB
GtOcx9uVpc/dhozocfhdj48BUfgYwG3kwcyXWXUgIxbOfY+AG/wjeRv0d/laq8e9
JCMv68/FElalB89QlIMYibafAqgEme16vrugeKFjPTux8kiJs8d3esdzWdh9wK4P
08S5KP0ZSMDPjTmf4EJBUEyh3etKMAccsjQIOhzpmDsx3ombsBi9Laymz01Uxf0n
qwQY/XN5Ms1f5PQHv8y4zW2VR43cWgJmwVR+wSWOBvCLgGlZTEIf4c5vjiBAfWqj
Nn7u1562QvotaHvLx2bcx65tW96wEvlL6nQuTKq2LANWXTye63OPghINdAQ2NaBJ
2fnpkmaofwLRX5vR5sLR8rzsw1JbS6TDV3y5e4IDDxICGWUy3fIJ4nQOiFeJChss
0EXYZFE1InFscsJOfOVDs3icwH8ZNW/l/0ZnQYY3QXpqWft2EMa6Ut56cKFEsghN
PfhLaEODI4bS/y+kwzlME5SPKtIPNCK2cS9oQiwU4zfxHcY8breW2II+geG9vBMF
wIJ7hhidw4OIDe2L9kLiKd5KcMNVuP376uWZYertrw45nAD3gRMMzqWQ5mb0Lujj
ORVTM8SUrAYE3Gw9MqK6eGNmUUHCvtyJYV1rU+q+qSk8QBA/levC4KzRY9bLxBR4
4T4JsMXAhpTNoYUlNBUzjeGI/oL3nD2OS+jzPoVjtJ1T5VS6vd07agIA4tdNxbm7
zbgc9+/JGaAobS0v+kM7EicXI4EY0aP3EwWhro7QN4or/Dthp82jsUPPQwLeQIDZ
kDTR2FZAXB4KfuXlayXmltBaln/MFVOoFcV2e94YJZE5cd4jmLhMSNW3W0KtUgBt
9AYaV6fzWyimWQ/Cn/1agyV/FOZowQUwriQkdu+lAh9WmdmRbQweNR4BoIMLTTWD
MzVeZGq1LTnnjOcJv6HirmprTtEMDsSIH2FtVdQi5ksOC4Fs/Seza6ufTbOUEudL
e08cHTdO1c6ZBeM7zcXfxc7bXCAm9ZWxQCMksr+TcbuGlKvqe+Yz5d6UPanvYAm/
1juYFDmCfwtwhFbCfmDCfgMXqhPohJbGLexRxKMF28OlJWX4djzJWugfHErOgB1b
MWIRHdoMzsB34KShwbW+LfzdH6Z7L9H5PzfqxGmdwgzUF5GECE2cbMeT2OMnfv36
4JeTfzHHyVwH3Q90Gr3hZKFoJH+J5DSF5E0wdEEH7rAReUHh4P75nueEA4p9rly/
rfHoc3tkFRioWXQJ+ERy2duzmlN8Zk2vPCR3+fuRqhzcqi4poN9ZcrjyhQ9iNMi8
8c36Lb5DPZeSVhSpNrB5Lol9TdhnCQEpDGI1sX3vmezIT3C1lMtgSCGW/d6S/eSR
z+UNqHWjyikfbjsGPeFpXxYeO4Jhxs1YYq5lEgxEqN2onachzEjpA5Nl/R6resRK
WdShUQONGT9z8ZlCVG7P+vI8kYUPBXPIvp4ivURb+fKtZtabXaIXVgk3vD8LbEoG
5TqukgEqwGsws4eEpACQAXi4iB768jsSe/ccB9m7M0NbB9VB9KZHQJI3hvQgUeFr
Xsu3q9tkd8gtdYSwRG/B5W/GRgUsig0SBYDwfkwiwaipW63iUUz03rNwuXtr4MD+
B6QVVdVjTuHoP4XLIjyS3TQWtvGeDHeLH9qbkg4azDYR6LB3JMd/hQSR8fcZXo0u
EtzKXItY7byoAfGm8vH76cProCy8o0zJUCreaHfGNxbD755uJuyNRIROXAalIXc0
jQSsScu9cd0tQ+ryUCE2/vvU0J/5b9uvUOFgKJmg3M8y7WcY7crjTuZr0p2J3IFv
DME69go/VLnKS1b+XSFR9XOfR9k+ia2MtEnWyJq+xP5a/uYguDP2X9h9M5S10Nqt
EyPyVPC+YLsbQ8dEbAKD/oKYKaR5SNeNz35nV7N4ilpXwkTcH4JKIV+KOBBbNVuY
0wQampuFpm+5Sg06HZ/aoy+HJ8mJNIPB2kgTV9W8+J4PKYR54wAzjuBzJKbiGyzd
Y8zNDR4UeVuNxy3G287CcOBqzHvtmA/RCEPIpdoPI1J7UVT6kCy/4K3qa8U9Nt6L
tjZ5HZHJW8l30dC62Q5zN0vYj4+xw2k2JVSQvhnnkx7MBUW1u0vdSXDuSPQjA96U
AZCnAXx/O6yIUHdLRN4lZqwe8Iqu6ojLPtdjICqMC+BXZvc1doeK23V4C3Sl01fS
P3aeNPnlKRdf7braD6c+oQ==
//pragma protect end_data_block
//pragma protect digest_block
x+Ka1C96wcbBtirECRjG0w4MUW4=
//pragma protect end_digest_block
//pragma protect end_protected
