//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
QeuVkIQit4H1V8ZBmExW4S7Cep16UTa+fC9tm7YJI6ksYIehwwtU+eKvUi8AhntG
X6jdhGAN7jG1j9uodzCkcCRcoNCjcvkSaXFlOcMmqSXYNdwPOnXAgWlYppjB9rSf
Hw8RVq1fU5BXr0ETEVcnSwe4tMSN1o1TWQReNOc767jNcHcBkdpBkC7kxffHpIeJ
HLEJWkjeL31RdRI7BEweWj+YSnu/SKHl17uS5gQdGQKrbOtwMVxG15uY9IGPLFIQ
Ifsz4daVHJIiH75Uq7kGJ5Ar8nkKqbGqRsxtoID4WZ4sl2IyIeOK+oC6wTTI66Mx
w/4H9WnoqxyWVGAvjGyj5Q==
//pragma protect end_key_block
//pragma protect digest_block
tcZE7nfW24TNTpy0aWFcEmGMrFU=
//pragma protect end_digest_block
//pragma protect data_block
pQJY9WtdePklarFs9KihSnuG3rg933cipuCOGMsRfrwzwohqsHMIgUmf74f28zZg
ybqrHZUPbMjaFpSQTZQ26baxc0PR4ced/V3EZLG3G/urllIDXHMmlWLWn9tMR3eS
rp8ZG0pSxeW4PWNFVTWZ3Ax+BH4c2obg5H+l14gOxh7UQpp60iY8VjtrqIXoIIEf
Htk3YSIFdOgSCD0np6vA5C2MhwHcyQp5aWNiyq+FLuwL6+yHEnjdfkRl++p8tN3E
dBT3IgFDoJcgVFNJYrxdM0+T/5d2uRu1pFUGITL+WT2KjNjGSic0a54GgLolX2tg
jPQz6HqE7ZY/C+niCgwXfQ==
//pragma protect end_data_block
//pragma protect digest_block
R//es+HzorqAp5VGZVl3ySjmtbY=
//pragma protect end_digest_block
//pragma protect end_protected
`include "Usertype_OS.sv"
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
NCRuUA1olF43+4tkQjo8MO/DBlgFDRo43pJQgvcxHt9nysP5BBAbZvlkM+c9B6jw
0dxdi4vjyGVACQIo7U2BkdhjLRAiI+Rq/ivSeHro1Lt2dURa3BtYW9QhujKpDfgK
scV04shSmaaJ+chSYMEeTmMKghIVXkSLdxPOfvSptUPMiv5Qr48qaMucbYRQdfJF
1jr4akraGJK9BFSb/Gg7rZR2yTc4Q90YEomhizC1rNFWAnrXt90z2nUqO/EbwdE5
Vys90wVoSC/Ohh4kbcp7/SEz6cRbJieuys/KVxsC562bhfyI9NQ/IUgF32hSCfNf
YxvUZtMtkij0XoWNk/JGSg==
//pragma protect end_key_block
//pragma protect digest_block
eAtFA6GhT1qn/L0v9ks+yDqzlAY=
//pragma protect end_digest_block
//pragma protect data_block
4XBeKCNMS3dTKoQjPE13p7VQUej3qmXdqzRTAYAVHNoxrWzXigHRbg01HmXResRB
fXF1nn3czn2GtQmC0clZ23mCHF92klZxwfuKskk4vbedIdsZ7G/BYu8QeFAQC9CH
CzLQ3dlSoyIo+n3dqjEwHkMwbqZeoia/dwIDjKhWuV/9IMv6UE+gFgrzNcFNsdyo
ZlMju1gk/XjOQqCyu18nwZ1z6usCksdP6yjtA6IIRQjtiExZ/oGsCMRaLdBAzozr
5pdF7hP7lVggIKXXg5VYQVy7YSzY4HPztTVJnoUgcQJxlDT+hXeOkw+M23AvuqF+
hnirnp/WKBMKDbRgwEKL+EqwqHioXZQqFP7Xb5UbL2CYZSFdpN/YNFRCMt8qW5rL
3lEGXqQC6wrmzOpXhhdtBxyrSjZ+pCCRhPz53pLLXlE/0jPalhlSPwWjBl3iSLwr
ZEPudEEn0fu49/6+fZEVgA==
//pragma protect end_data_block
//pragma protect digest_block
qTd/PJsxe5cU99B8KrzFsJ96jEI=
//pragma protect end_digest_block
//pragma protect end_protected
