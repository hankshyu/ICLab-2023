//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
d9w+yjRAgCBZDejsC3k8K63zqCg1ezn280QY6Uji19ZAXOtgYssB7Jm97g0Fvua8
FqvDqWyRD4dqJCuWcWOm4AnTFTgVT9oTvqt7goh9eMAMehKkPNXnzDu8p7m+If6a
tB/EXiS8OHxnFhE33emNsCfNl5winN3KkugxAuvtkUTtN08AKDeRN9iqJCLKsh9G
RpEzc8i0ojs+RAK6QCdoht7WVXkD4d0GK+0WWbkmaHA8zBtN/NC2T91KhMZe1gNg
F8ndM+Ha0aFi5vwrbAsJo4SVQUhLHuEt6SYhiwqicKqPhx3Y31b6kh2R5iG0Z+El
GN00yTw6ttUKB3NHXXwkkA==
//pragma protect end_key_block
//pragma protect digest_block
h/Vg1/hbyOYX2BA6EvtlkDYm30s=
//pragma protect end_digest_block
//pragma protect data_block
fMbyUeqGm6i+0adgzWbq7eEDnnf2pi5niO2h2fC70ELBs7y6NaWo5AGTTDDXWsRZ
2wdhQtVleLLKqRHD7im6uhZdHeyTuoQ8cAjmBMUaIGj+v3WgVvTGQ8szn4OHL54C
02PA1O/DZXLJh4e62Nzk1dUdPiJnq1CRKb2RD7cee17WYfXZYoD8s2yi2BPH5qeL
fI25r1IyBTjPiGWnlapXYsKeJLTfci7gVc/eZEqqesFmyJ0xEjMTqjYREkXgf/WQ
9IWSsopwCeTvNI+DhUZ2c1219ayOOPbMooMjuLknMHRKGSDoQOosMexRoDqgq/VK
/m6CqBLvi6xC6MpUu6YzMQ==
//pragma protect end_data_block
//pragma protect digest_block
utwSGFKsyEdFhKsKvAXFD/9cm50=
//pragma protect end_digest_block
//pragma protect end_protected
`include "Usertype_OS.sv"
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
hmKuuwPAsTcHvpqYtPtb0bAnUo6/JRYLa/ZOPRuF1+tLzmbRoLTfHe+r+P/3UZWN
kl9pm5xI4kmzV4s5zugWd8zJocGgFBawK01MG3igjDKmmIpjp9iY/R8xg382FHfV
YAzT9jCNsAsWuUgS3RhS8DInO/lJV0asaZyESdVmyLqxyjrCS04bqDLWADa/+0al
CiBGwok4r9xD0K/VHYO8Evyj7FXFkf+3hPCkKIIQN1RDqhZ6FWGGwZ9lvQE3t2jC
AcnTWgb3+WBv53BzV/EFW+OUgS8yVzj5q6kToeij7g8lFcaUrtwUW/JYWFw+r6lh
v7XHkxxm41krPOzVrhleyw==
//pragma protect end_key_block
//pragma protect digest_block
2hOnhIkC3qn3We5Pa+MlSrNPBO4=
//pragma protect end_digest_block
//pragma protect data_block
npGvL0++e3XNN+2Xv9vNojAgImeEqyRpIm9iD8VC4p+Rgjp4KLaHrujuHnAx4DKn
ITLuOb9GO1UvEKLAo5ZEpzB65Hr0rfa/1pWZTIQdHAniE3CcrcaGm3nqid7Okevu
LyrHO9XpZfNaCiSIrQuKhZffHcqriG9hcZCJQ4tqF2XbCJ5XmTo6OQpk9EVvm83A
W6Ugo6qEwerjva0Rof7F8Rjpmj+tuNCnbvOaV50z0GKU8BXdEBnuhS/odZQXGkoW
JuHmYQK4oNCRufJsRF6n7T9fFOyztSL90xHkpK1t+MKRtrLP2oOTQNSDOn/XksPH
u7qHyWkM7nTehusHvC8aRETsdyoS67Skc+k657/OUDk0LsagggLN7oT8pLfAbuBT
TSH170iXyb1wClL/+MyePqXN3S4UaLZmScEzvV5ZyUh8q0QWfnwic7LUigxBj+pt
NNyUNzE29qrHI6EEdzolf4CXVikVK9/7jV9YsCUP5U4++6rcpHixnZMEHcqGRBhP
fCTr7xvPeJ4No37U+22zH6MrMgyGtNxuf6+EtTF3QGJZ/lmsIlNqoiTlZ5Ulooaw
ka0250bJZ8T41DxXrlFkWgAmWj3fqM9xtwdhiiug49SlIxzqlFWXLsCbsZdnWG3x
UFmRNheWHaYYzWXaW6RgojB/k4BYSAWjg5fKGd7oNg5XDYpRIaYtLIQP7ynVf8cl
cIM2XcS99/I+PxxxDM4QzI181KYmxjTn7zMjKWXBHW7oGFW9PAfv5XH4lUoJtnnZ
2EdRfKkhdJacugO0ANxbzq21IZ1e/Xwpfe/2ltxLsuEdPdGqGxi0X7DBvmpkOo5V
VI33dlKAAdoI7LNrY6uN2/YqP6a91z3wA4rAruZIFbU+Wkf4soq5vncG3sVERgAA
scUVOQwkSADDOeZRfKFDC/30+gGgyjhhcaBQFZ0Q3L8mE/pccm7qXUprLGBRrbod
1WEXZ7sJfXdgAA0TavQdRoM3zYqGc4UuQ4RZuBeNXyy6j/1jKFccvtkt20VpuScr
uHpcoJw41OL8rAcYH+dABAbF/TrJWpn1GWZrcggMrdux3CS0sJrMUnOzVR6tACto
Pu9TDS5mBRt4YlZSnxd53soXoSio27zVDyQgBiKJEL+OhG/mhs/gnN1fIdxiQ0F0
Y9YmFOEQc0+0HGxJt/YHCigoXr7a8zWdkvZ/R6HojqM5Hln9U0AURG69dvkkDLeK
Y5yMr0hN09uO3EVxqnC9ATz5glK5UJaf9gbRzffmkz/tgufOol23iNerUfh/0I3c
WdZmL6VLNM+etz+GhcBEVJfXAaU1VE4SglJnQGai+OIiyj4m4MAoaSVQxSXPgsrZ
iG26YjC7MloAFh4olkG0IUfZmpAidemvOQDg6IKuvFkRuAoD9SpzuaxQT3vjvZRR
gOq+7TUyoZN35IhPmzgM3mRGZYtOf3RBgJNDjBdTMUAP6kPP27Y56DqzI/Z08DfO
EGoSMtnSwDVib1m+0sK2Ec+CtDvD6ChjEofDx7WMs/ulMMYHjNV/UeKMxMfOCqk3
8FW6afx7c7NQ6xN27mHn0YbOPyemuiisUDIy4TuwUC64hbmHFsEbWVhcYCbPkEtM
PdONEalkl3GW66UERYO5KvIBl+aQBXhi4OJ7NEkV6GS54Bam4L1zXNCKw7OKT3qT
AikkyNbKlWn554jvGTQUHkEf/vJEWwTYrdSZP8UiMGeeke8Fqhao1g99XMR2smp4
CK/p09sHYGEG+HMsLQJtEWNOAZW2xa4ZwIV4zvvWnPcN39jilrmOPRJrGgtU/y8B
1Sd9RWLin8giL3/B9AvHGbKQcS1yT+UMXD5QfkdqCawYVe2A19/6ruSoHzYnGN6t
IOdXRpKOV87RznbTKyu9q+cFwSvayUqscn0vd6rPFjZ6sPU1OFP9MurJiz1Sl+1c
EC+VNZF1Cv8PDnz/tBF56Rr2KpWyld7vBWCnIZnzNTro7XTSc0RJ1zmLO64aEHPg
KSNWQIg7mEK4GqwpPcafx9YZ1GRvxJa53aPGoAtvdRibw15/8R+g5FWocHi+4Njs
oMTxvngMRCk/KWOxaxk5MVn3GV2/6/RkOinm/lqNrpTRy7CYnCcRELeFjdZwXR3p
d/GzanhebiwdA4/IgY6DLaJp3psfjgQ8ajtjzlpHlHALsIvnuYKXRhFeCONiWAfR
qzz/T9IcFe1fO6vK5hA7tH62XzVOuAPxNFVevs7gMsp+Y1KkTw2oa9gFZ2L0YnS2
5VFRgnD1EQ8t6t2AT8KPszCmeR2WwwTChhnUwdejMrvj8r0kRb9U/AOFW7yvekKA
SCdzO9PmMioDaGshB/+Z+8rubDyskcFtKkY1jRy3SBjox9c7QrnX5YyG+egJqX5V
IbXwskNaBymgdtiZ+N+SHfcYx/GMbG/g2XFO/KqUUu69iVQTUEWLPI4pIy0/vmno
zO5AMrwyeWD7VLXU23RbougigrfCLcuy6MgIP+j6eEOpKzdg+HNV2RYJDsiHq2Ry
Qq0i6x8skRxFIp5uUMCJFqDuCNU/KKdFF07fg+LFLNLliokRvqUqej9hykjiW40V
4jfEK7ae2MivG7PmJxO1Gw==
//pragma protect end_data_block
//pragma protect digest_block
vrKDK+Tl9cA/t2l7s7QCgpnnL4Y=
//pragma protect end_digest_block
//pragma protect end_protected
