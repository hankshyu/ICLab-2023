//############################################################################
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//   (C) Copyright Optimum Application-Specific Integrated System Laboratory
//   All Right Reserved
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   ICLAB 2023 Spring
//   Lab09  : Online Shopping Platform Simulation
//   Author : Zhi-Ting Dong (yjdzt918.ee11@nycu.edu.tw)
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   File Name   : PATTERN.sv
//   Module Name : PATTERN
//   Release version : V1.0 (Release Date: 2023-04)
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//############################################################################
`include "../00_TESTBED/pseudo_DRAM.sv"
`include "Usertype_OS.sv"

program automatic PATTERN(input clk, INF.PATTERN inf);
import usertype::*;

//================================================================
// parameters & integer
//================================================================
parameter DRAM_p_r = "../00_TESTBED/DRAM/dram.dat";
parameter IDNUM   = 256;
integer	Pat_num = 50000;

//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
fZmI+ogzhQlddGr9IZ/J2UYSWW7YVqbFlmBkwosYDy7r3bZ5WhAh0cnDxmMq10PH
3bnQzQ/wWhTFWGiTKkt/REMggDt9HmxJ7lmYiTcGJKNQ+RBN8vSODqtYXFBAovTQ
xqitLYmyPHg9jmZGWMT8LHhH6LS2GJi+MIzF0zCkUUPZquS2BGJzmBZkMEDAMvgd
ZlRCALnEvDG7NkRFI8V6q/zXSZDeIfSvuZEoS3t1ddD+BaDqgFMN+fUxab/00gNa
XdfnFPSRV6id0Mtir/m/vuTdketq5MOVZcShVLCWJGoabTg7k9mFPA5D1FghIeaH
oH6WhVAultmcUYPtO78ang==
//pragma protect end_key_block
//pragma protect digest_block
VYsALtpLMJigMzgAE3aR+8ML5gA=
//pragma protect end_digest_block
//pragma protect data_block
2+87OxMPQFFYm1L5QIiZ8JL5t88qsoT0+d4qYwf5Cl78jlEQ9Ha3pfEJkDfA1Ykj
/iu3lqTLBqi1hvn/1nQl0HzNaeqvkw2rTtRDhGAVM5YuQpR7EgsKhx++Eh9sBtpE
k5BGw8zlpptrUHIc9PVPsJX387RflCpCxmNRIu2t+IpqmEmIm77r1eb8/nMf+ReA
gyxfZ8CMLtTNlmPcZyfQGW1nMiCApeRHDhf8RXpwkfCadu4xvL0DDQV+G280/R7F
U6QriY0zpiwXgCptQA3XTKxz/1tte1tJRRA0JFae20NsxZGGxIDDeQKZI0e70K0D
dC2wG6hMckZRfNHqPDhVVWuYvGSGgzcTzvrnP187YU8cwzUuHf7wFBLqjEGG5OTO
mpY9avYT7zO8Dq+6+MT0UJhUDc4Wx57Apji8DwDnioAf95+0mwsZSNWPjz4BwK4k
uj6v/qkr0R4PwdHVOlTskcm60o7ak2m0hGimTfZJ/R+/Otv6kABnnTBWcaFjLxuX
/qKyEzsmnZqKJ2jXBP6GRpCddeqj0DoreH74C7wgXoIALvRZsLdsQIj/sJboGaY6
7GP2lL292WOelGWjv61zeywFJIkK5OjBMIevcOi5W4BKWLbTiLdKnDbsvk0bikup
YEDob2p7IaXEZE1Gsmgin8PxGCn/UX5Bz8MJWeHtyTNK3jR6cyPp1jUW5g0TBjux
VXdEVJBrxADibXHumAV3kDAhcQwp8v44FvxcOmnc7ITAIzzRZ4duVPpC1/wL/7SR
j0HyUUGoE9FJNLHFcXJFwio3XB5k4wtfyyRbDz395SaMXn40fEJVZgfd+G6l44Nm
yhPVL/sci2igfxL5akmkg3g0ZT8/2qC5f4UMlVmbMawaF1VpW6JwTluZ2UMQNasQ
uBtmBaW46lHQVJB3sxFiGSaUX5K4rsx0ZO1uKOyScCOgJIlcM3Xj437X1BZPfXib
kG4n8+YV2HNNzVJ8GRomDxESdx4SoebtdG02dvHIC0tdVIyit7+Yd6bCgnV2K+Kg
PLwvl7Xw0wkRRUbtawenlKxdnkXWBDReLxvhyXZHleAR73p7zeAJRW6Z9dpmLj8x
ugyJMgMzqkjmJWJ3goPVSmsReLDJtgYvrsyeuAq4dKGjomT8obXJKiB3Ax6byKCI
d70HeQZaR5WLdP4738seoQVIdFMpxWg2lL3lkwU3KFNg+Wl7Xp24sABAVifVUruj
maBiPwbCoCf0hnZSw0wtH6zlVMYw1uG4AMY6PLfMhWoU2zCGsTl2fgwRXrTXyrzt
66Lxhw14X6TljZbt6/C4lC2SLv0sqJ8aDErE2Mn7OoNxtOIUPF+fGKso0EN/I3i9
dFpxBxy7VscbHNOl+6OcY3N++VNOZ8winebNTtVXKV5sMvQuvHRu1ucazRbwAxp3
vdrSEBk8IQyEBrhTltCOs5dyOJzpA0GaquaqFoW4A1CzNuevjGH63RBpEH6yAPHo
qz+mF/Bq8eLh3q0jphnCjJE3gAzz0T7xbhMXVkAeyBC6F2FW5rocJuivnG2DLJ7p
cxXfAHwKS5+gEOUL0R88Rnulv2H6H59zjOsNeKbUu1lBQMh6sgi9V+U4dpofX79t
F0RcjH2wMdrNUry74d4PTpV4iRxGrXlGwiA1djvnS7PMyRbPOXDH0F2NLxx+ne9V
m6MmC5xNA/okxxiLR4dawsI0dffcq2ofBfksQ4dV1zf28G0TPj7De85JEqoMZFyQ
x37BpgBB9qMoC1uvinOEUpzVd/peq8Qzwa7usAmytvnb6GUN7Z8O8yvLnRl5Hdgy
+n3tumb707Lr4HVZFKCqJdKmFn7x+LGnZ65+SSmp/GjgD8SeTCswJgkMKFQHaRuA
y8kIVFs3Z118qaQXsNPQEPU5gK9MoSSmK9yhBMpkn73gyAuvOI3M5DCl8f4iftoa
Su7n4sTcfcCF5P97qcWvnQIAcU2Xb/8opOz19NHjVcHozAZ+9PyXbK5YNP6gziSa
GXbIFxORB80XM11UMQCAlw5k9hEoHiWxipxuH/PgNNC1E1Dd0u3E2uoqR4f7t4x8
yHo3D7pVFStuyoq0SyjLBd/p98yd3s/kwGo4BS6nTVU+mEBolMpZ5A/zNZA8pAjq
zWJSNdR3T0AccBnfz7MYJZq4ZX4JzJLHqby+CTE99HZP+4qAHKkKR0rqBy+1Aboa
Q5HNA9Ywrm+bq+2n+dYI7HfjacprhITcP74Hd7MNNqSYhJbhxNx4FIPz4iAnBP6R
rI3aW63msYb8fWsPu0p9BaXPyosCgeIDbKOxcfBTvNgr8WCRXXoSYl7mq/lrRGmv
lMWjDK5M/nilmiJ0zhq8/x/7nc76q8LVo2sFvVRUPLlrs+X6WBxnW1KucHuMo5Yv
O1piYRpUtjQTRmR/bSz9+Svr0kGEybS6yHFOyAZE9mkho5/Lww5WMacqJlatDj1M
7MTVB30sTfC/5x5AnQbna7ND8JHxfpL9MwAGHwNuI+/FrIDv2XvHH7UGa4r/pp3u
A0h6xg5wOCoC7YmOW68a9SfX5Zp8HKW6pqL7EfzysDDZb5pcSKsDQKIE2txAXcqR
OcusqWFJnMet1Zpan43eySzfmNtnwaWDJuSqce3dTj6sbDKfdgnOmsmHQCF93dfs
bbUYT10FLt3asOIZz2qPQYaLg8lD+C1fjA/M6GkjPNJl/vtV8hpBjSIvWTNiInR/
gjiQoWYHaMq/PCXUbKcx4G0HC5vZm+s6TkweI/bRa0JHnNHQuB4SWmJFGHSRXWN/
RL8uEKdxLoZA7GH/mO3hLnbKDBZOchjD6e1qFn+BhddhK4iEnM2AGK6z6nzWS3OT
Huc1x7nbXrtjtjOz9c+U3g1kTrlRFX02Qignpw9KcLGAx0L5Vnh0v1mAT78EJ8vR
mbIi7UCoszuW9zBaXZugdoh1NSm+NYY6a2i+bux8C47yJfBWV4kWo6DzLSME43KI
9xr/VR6RiiNCb8vYgl1jPx0BISlLJ+L9rma3DVts3M/ryHFL2lwgfFXG1yeO6RUI
HBGttqPR9hQhkz96r0wEOrg9Jl46HYpATcR+Q/1YWsLcJKPAgRFdpjDyW1Wd4koW
z6fSatIJlH4oXp2rZtKhALPspEPQ6sJ9LHOIfmZ1SZWS7VnJ+KYgooibidRayLmp
xv2E6Jq8qcwfslEiuUG1EioyEYer/FMPe85nZeqyOaBcVFlhGuKEEhqrC/wsKwwB
6O3zU2k0q5RNDJWaggivCp+dhG6zxtfKgs8QdAnV9aa1GAx1inFud54cL4jY/wDG
rYRcWpvPNfzR0ODsSn5zoJgz1brNiNPwPy6tWD/3C/h19gXVobR8wiqz6zBUsxPB
uMTo2PyZ00JJvDJ9kU2DgCaI1fKLxwQ6AG8zsBhoDkXy0KOM3pYqE36UUQRVnkfJ
tXMQdWrtYGxomGOypHEiEkKmuSM1ksSKiwaYh4tfqjtc3ck3aCcFrXO7f51i9JRS
XR1gKgpVFBA7Z6N9GaST6EEi2XSOeumcb5TRnb0m2enRiERKihxFTO2ti1gjYjG1
dVtY/IGhGrGvC8/6IsgH/O0xyhtZWHW1RGFo266eDxktBCI1nN5aG9llILJC6xCU
nhyJcup6tvRDTkZ6b2wuHqBcaClHnvwJ3rR7+xij7U/lcHyEyxc4uPhPEvu0j/ba
3l3Hbcda2TfQclwnmihKipj0kupFV5c7QMQtG9JcaJkC9ffJ5PQIESsthHHHTVHI
kmYkBmTF7E5eCrXJDlTxBabBKbxds2Na7tyr5sj58LrkI5Z4YyvPrvs2y02I8LAI
JIhbDZrkVJjqARF2i7xWvmBXt76/NmUEH+6hSiNeK4u+uAGSx11lwiRQ6vPuz8ao
Jb3q8Vim+/GPtiHhNdXVcl0V8MZ6p+RBMucIPK5sE2lpsbmhSsAPmbIqLQ1qfJll
bY3lDi5GBrTTLdeA01uEHm3fo/OpksFZo/fbjBSL6CjiyX5wLLzIYG72CddMajwi
LOmt8XbkHSLropMh9t1msYkX4pehZIFuvlmbBkX2ktN2YQwAlXNhzvMUTUZ4F3Fo
funbi7hRAIFKprG4zThAkdJ5UiAFOLFQtuFjCiA7ahhNmQWgWm/bxL7wQyWBKHRb
v1aVjeba7uOSTDDMPCGgJ5ubqmGOE6i5XWH3ZT7jG+XXQ+kYL0oo/GWb1KBoSXva
nvIPdvEigYBHFEqTNqgYxZaZx/qz74tcDlbEDv2/BUmtmSxGpWI79V5h5T76RLtl
CaPF49K32QYR6teH5GgdRpMWTg0khe8cCytyGfOECWTYksH9RolO/TrA2ZanYrE0
1OXqcxM7cM8UUR+j+vpshP/TN1lomDwgnk6SERho2bpS7+nI1Y0b5GJNyFollxul
I/GtQqZReESeHSbs97X1vLIi/XQ0dQf3QAqSMtrJS9vKMBxppqEfjF4+VzUNen2G
iC93iMPPfHmkC1wZJJXSLywyffGdB0G0XijY6nyYMxOO9CCdrlKQeYJoZFhkaE+e
szueGZ8E0nNk+a20DNu2o7n/8luV4nMoI8S7egIavCa2b8HSuZebOArm/TrMm3HV
3KVoifHvijYGy07EsAYTR65rE++CKSF0DNI4LafqWo1J4THF4wTJP1hZjP+U99Cg
DLeqyqH+LNhhN8JZbUfHna4ZmczoTeKj+KFTolsjUy04Ps3EZfhyznfqWaCxter1
HtchFiDtfhYPMn8KgDvYHFL2RbDEkjCyNtcS0gaIWu3ZS7gh4R9FhxKEgJOcYn2G
//Ng85T9J7H7GPddLCLsqJcd0h8VxDpvoIvuqk/hJi27Q3KZXC4nBhdpp5D3gHLw
AlYxigR3fXWBmH6TpCg9vo7k16/YSL3PLguJzuwkQU3vYAEHyTvBLKUUu94sXNUx
k65bd5fXyZQkzEN9JAX/JwEulPf3g26zY1pcBoy9+OEJ/soaGk+0GqW8g/zLlU3w
ue/lvDYw5QQ1s5umvst0xXks7N/A3XzIXmpt6IwLMiLw63FrKPGmf9ONErLvxK1P
egjmKv5ncC2fy11ojLTJnsqnk9yOu9l6Hxk1LDPqXlSUa/0OyIXlVmXG1AIMWx4c
rrQXtLguovPHppCk/yISJvzWiOx9UOgrVuCU4/WVV5W76G7SNEsLMMrIZ9a67nnu
uVbabSXjeO0Y54RbmDbfdGWGgQ/OlnI51Nipa1nZY28ERDV4SyjGooCVhIQkvOfq
+Rc4Fdnasx3rqqN5ErReWAYtXUv0C6nCa/OJq3bfww73Yi7fPVm6ma7LW/tQFVQ+
1lNm85G1isZGIxZdEKbPCmv4lY6d9Yg9Iql8sPuwj+bV2FPSftQyMZo5hs4PJTod
J7JgikDDQ2tpCsVUKD1kMnE6vg6iAbK12ygFcRITIesrSVYxwRA2RRPb4ZsPB/hk
He0Ko7BxwX8U30wFhYV7Rv8UOaa20NfsxNaW01uSa334qQYvNaTmcJ5nRg3wrOMR
is8s15fosvVxFT/7UDJ8KYlxNlO3QSmqnjkZrZz9+M1SCRPQ6BWi5NcCwoTuoeQT
etahphMNp+Q8XEkHq2mucURVLDtSiHjyZc9B69s4FiCakDO06CtxlQDLATxnlnLx
6X9AWt1KNiqofKzcqK/B5+B+l2p8fbmi7P+PmLdpW5f5y++SjoNmmhgLrG56HO9r
eskW23csYy285MsSGRGBvBpqPdpjCAsYhziQ11SLDVSz31UAXg05cp3ou2Sc6JaS
x0dpDfsfwzBfN1c30/ksQFD26m+qegleoWnu1g3nN0Lxd1++E+ceGZllaKnf6PTB
rgXoRco67igTVkv/fJTOY4hhPTDDQnCM0ub5osmdRalLW+GcB0KLMvj7ZmcCZtEd
iTD4ilXceQWzluYYt7o23GmmXjxCIRDiyYgIILPTpQiZZU4Rk+WxmyTJY6GExD6G
3f2C8419QbI66gsPjbtZLmiSytqV4tMDoDGPwPsQMxnhkk2pOb3afj2sieVu58Jh
0wAiuD8mwYDkH7UwLfELe59cO7kit1EisckjHLferQlbVDO+v6nzdbNrz4tK9em3
gEaE6d52UtN17ubTj/uB8f7/amXiMODt8lHWpIpKOHec9mdeZUelfA2xNJQ3tlYl
FGQRYxhspqrgevR6zYTxOttruRfuiMcH17h4SIxaMEB/YDaS/12HhmjFVtKHmi96
VaOkcA0CpRRdKOTkXZHHK7vB5gLbEbM/C/bfh1aI8ATsgAXPEKrfjnAFGb+pseTk
XD/O8OJOmoGmsye/v85qzRfafJzopvNT1ovqj9V5KhiUuepgmnCnUgnZuP7vWTag
DM+Fn2rZD6AOwJQujK6HD/ndk+pqEYpcjXvJxc65Rmy9pFXB8W4xXirCJ6SJOiSC
kxpt1sPP7uGpn2nZd7dnISfcud9jcjADH7V7yT+7Hrg7X+q4KW+qiZ3xTzyK4Iww
e0XzIwBbytelX5mqaOG/ImTy+MSZv6xg0p5Ke1c3hSIcwJLSqMyVYW+BgAJtt2s2
dzhAk9vyrN93YwwEPKyTVwnUTgc+XMgCOHkIcHs+TZ/+zOFzlb/k2dwOc4u1BqTr
gNfjjny/Edg/FTwMrXll1Hw2guEbp2jZfqbR/bFwBd9iyCTuN8RzVqdLwd6RLcP6
Vy6rNyyyjB8QImivst9IKNgDHs7N7GqGMOjezqbpmalGW9mqgzeCkdm/0mKg7wPz
VFkLwtakbwi+vERLd8kK4WWniWDP7mhhb6HMrxLHawzFvAHjIVXWumaf9pUt6syX
2pcv91Ej69E4opOZ2zL52U06XHzVpxbCpamD9KPjAiszUUyhLUMy+WzQN4hFJcvW
9eZ9P0hBwBY1wfbBKkBkjoYET7UjS0PK4X5MhTVDH4J9ehUCLCAN7FrVrmHVmKvQ
DbaP5LjuA/T7CXssgpPwW8W46F5smauv2xX5H6JO52hXtzD05C4kV3X6uFtssoBi
5Iybf1Hr4jVUVY36cWpr8eL2C18y8oAe7tOOJRzIY7TwunnJP8brf94/0DpHDAF4
znqx/9bAWRSN4ubSbEVSU0N38OxC5qa5cuX/m9vVSIUmjqBWFr84KOjXjTVn5a80
8K7OXsTLWM0TWqillDZ5MgLmXfjnQi5RsC60lWOKy756rhIDIL8NeUTJSwyBlw/P
3owCXWTs2FtNqPMU/ADS7O7bBE/tDtETdMAYxNS8zEbItm89lFJZoLTGqES84v2c
mDsbLsYYk19DbbuJmMrVqgVK9vd9pSh1qZwqrCX0+IawlWy5cG81UsFZ/e3s1Z9i
NPIylV8j6ocob1Z+Z+30nELGrlZ18inyUmhqsYnHuWhpD2mKCVTJBJpw+uuqtCfi
bQZYf4larl8niM7xgpz0w44aJl0noYRU1zz26sB3pouD+yq/Q69jSm/JIrEYFvkh
tHL3fKdffloJKYaH8ARbiNnw+0mbkkTBnTVyt0tRR2H1hfTHgDN0eN90POuoXGTq
5TYYTlExjxGpBWGcyt30Y/Ld4vuHhts9a7s1OuHW/pPZFPAUYGDQ35yy9QKarhL5
y8uKzmnnb05mop1toka+AWv/Q5OkHUCPk8ZW6TRV9fzB/h/BU63aYfubj8DgOs4a
N+DiLsy0OgS5w7WPg0f5yL5dG7ZwXJ/ENYi0D2RiljIUhnog6D180xCMkM2JMSqP
dl8e7GC4fXukJJZfFkYjRV39ldaxXPxcQGhgZlj3vBn90bFakHpdV0ll3DptiOr4
Y7d6D5ZOWpWO1ohrMYx889eDirnUULWtFx8XKprmVwxoxDQVxeeAfq0Rw5H2s3Wb
tsrJ8TCrura4ZT480OJb1J2XHmErqLcrfcptIvj3BOnfG+SHn5iQJ0a2vKi+/tzs
1ZEIGAaaCzIIxNGp455tYSiPwUJhhqxb6pn2WTrYlAe+7Za0G/gL7OhW44qK0MEK
wFO5Mcrp4mjWnyCfMm2BV2nLS3AP/TnO6hAHiyFiXcdOZltQv6YLlIIalgdA+Lpr
AP45w/JCAfOLXHAWFXGrKc1lyF+Y2gyMmu1ZbqN6Rt4RKJPxvnCNLo8SKBOa7wfz
MicGR/fU9Zp/nwtZZdIBISaQs4+Hp4LHu9PB6+SntUgnhG8fJ/cVuLEk7bgDi4lU
QAzUQQfkHA3TRvA6Cv+8CXimm9zSmV5IC4MwPXa6NW2IXBOuuV8Y+AOO9MHU7stL
JGcGQ4ESCsc6Tk5tEk7mWl772uxzFzPF7u3dy8u8ihOplKPHQtZnr2o3eMtzVF96
qU0SPNBAzBgqFtb6RtTN9KS0HMGGMZ8kP8CKiucjdLYZvrubMPLE5xj+L+OwoV5G
HoKaUFDnnx7i21MfbVqcUedMN1dES7wgrVhZIJZtP8LgysXvGiI4phZiQ3t0vPjK
b38mQV3z8ExyehWRzNvHE3kXK3yFQEfPWFtQk7ZLukV7CJf+wcbJAvWhu5ZAq7bI
0cnvJ8r7HWXMPjFuY3b1SqH8jMqxCF5VOXDO7haes8ikgL62j7nptQ4g7Fj669va
ys/iubVa5WpmAWRYQkj/0Yc61N1wucDa6VBo4wgrB0sq2LFM+v1UNE3dxwf/49CO
41vTInc9a9CZhYReJKNg4XBmdAF5w+hU52IkG/r+ItA1bzmUa2PgbUaLyp+QYgVn
jOSOJ5aFxOORalf92TqbGVRrDrhjoje7rKMVJ6tKExUEGb9oRmc71/Qjqw2rFu3B
0aru6JbUnx32+wEfCKprmE+PKSNDh5YJb8ykXll/lDpZu1cvSwkfKWjCexlUx/L1
E8orjqEPWY8Hf8qSoY+oW365syyyq9tDbEczoRXDFLQXyMKd3Q503fPBnrVUx7bb
QUAdDipyRS9A3Sv29D0Czc9BjmFPZYIcZapbGcqXNwWiuCs5WGut2lwWzQ01nnMg
tlZX/Emj7UpV27u4IllS+AGshK7AXkhgXEfvDrxeK7nacM4Gu8av8a7kPVIY2xCe
YPrHteMjj+aFjgvUefyXHsY9kkbSqdSLgWRz37Ng35v0E5xnQti0ZTskRg5uCDla
nNNZNN1wzNNVSlBLKmBJESHpPFvrwV46VGE+NSi+yx64q0KwjNCdqHT2IJ3CNVK2
wha50tZxsO5fGA2lfXmF35RjJVrl7/GTOZcMaRG7o6b/OzKkLrFf5vob8GYihmkz
J+X+AYgPgnS7GZVPDDBwkxc/JKUO/ARVVhkmAnhYSYsgWUY0DYBsxj7wXAxBOWqb
9ePx7ia8qTJ0jEwUZVtYZBqk0s5ZWxHxiSAF5UdVCXE7bJNIJ4aL9gzEtvb3irsQ
dVSsdvjU1tu2N8426KP5V27A5Kil01mg3ByvblvIO2RY/jPwQ8Pg5N1QzMI/s8nH
kV98fHmhZvfi4Np/PwreOfBaZ+VNbTf0dLhzllRVRYWCn51dRfpRrPr44MKLFscF
pnkh1b4Hz6gQvz58BgPgW6KgjuUnTaXgxlHDAnlZe73iAc5IfA/lkOxrS/aFoK++
JveyeQqhhw2acXracdOHODbNsTmkEgJZLu2lwG3wx7TIH1pr7shjwRb9sta2O3QE
SM5YNR8fK6qHttHF5CtV/gkCFjKb/yIZbj7l5GTJX+Hfom4tg8oVMFe1Lg06Gdo7
fagSC54O6jR5o5UDj9OW7naxRXRoS+wpXx83XsloLXo2gOB9ervB6PIKNohKOrKp
iIY8K0XuR736s5mQFqqNdl4AtxqZZeXVvrfMQnEbEWzuGp7pFVT4PmEIR3vc23d3
tUkAsWeMWT2d4rRhjMOp7l1+MmX7/hmknaE11q6ecrJ1PFYChBqF0mJAdejXltjz
RyVzAZEHL+ZFExNFycA360TwfrbEl3c1fSWxRwUcXzq33MY/bqbf9kCECPn7WN4R
NlMqR2L9hueH5C/ra6gcZFud8p36BRUKKPgM7Azk4pBLd8EyhjZ+kNClo/UmZsLg
a0VLXHVBbws/fL1HDkLkTGn2wknvaFLOBw6rUBreinfrN185UHqgXTve2aIVp5kg
A5jREB/yKyKLnQ9yzStsANYvVfDBTudSCUBVD4H0vF28xaPownDNQEPwGWJTJqco
zj2D7tKYI8KTyVLyR6J63TT79gbf/eqa/0gn0dI9AxNPpacEcRZgAMKeyTieKriM
r3fg88ZLEcni3BiTlxrU7+1Rohd4qI3irxpn9fFfY2446OnLp2EGEQPbJFiP1zWx
QDGTtD24wrCV9lwbG9LYnkezlfDMu0Sjzy+AOCnkQIpPHWXvSHhJSylywB7ZdQUn
Zl2fQVK1Gul6MFXFW/UpGz1ImiGSuXbVooh+J9fN8F3JHHBj9sIpDP+oqRweDN1e
rTlzdfvcvB0vSLhuXjgp0cBNINBcdw+nb9UQyGraifd4EVkZ6WO31GXQ6vSHYwy2
vfCqeKir1Z83DOVXCR77R1kEMFdMjcEbmspjgtQVEsx2+SZ8YDsC2gMIrmHrcTBe
LO/f6RRg+m3DsDAiohWK36jHomeRthDWmR0IfjnwT7DlpBc1yCgVLeUpcohjY11n
H+eraNIPKKHITTy41HaJy8nHKWKlehyGhzmaGaeUn5QbSyJefJMySahFaiPAw1mV
YAr7pOqBL1BlsDe0MossmDV6TR44ZUujrMdYQ3HnGYZa9mqGcaPKYuYsoK5VX1Os
brZ/W/4TlBk+iVC6mGB9R40gLJrWuZ2QVAwuAfebsWowG4pX0nrfiry1at9bNVmo
SqRwzKMk30oRTPBlpCjXNAzxmJPYXUY1Oa3O8mITzLupUs/XyHWiYHC58UIKdljb
x4paDlb6l65VDtrEPM2HRY8ACTVAMXmJYZWqOU42hSp/OCtZWbatUDpjMetQYFhx
u9vUOaxDB4xhIvSbKUcuTQv66SfHtr6+l7EuFwXQxahq+NRPi7rWhXlnbfxUrBhD
TfqtYyL2LpVKOvuo+ZQkn8BudA/tlARZAboYyxRlYRSWezFZNDnSZVcKfUMQIhwF
fZzUJRpCj47iqaAmT5IJuSlF91D2VbU7JLBa8fz+MU147CTXTDE1G8w4PbiLZ5TC
/Uc52S8kaknZhERUvvEd4wz7nm+sXRyyci8knbuNiNVAo+Q3evEoj82aOOgNULvz
o2trgTiWYhQqEvZLDN1SKXPA4iBEUAF5xN5VzF4DKvuoG8axY+b/V6CWsxdUw0nl
ni0iC03Hp3UscsvTZGFHAbK/u8a91nAhfBssm8nAA3HjJGFKCMxu9Ls7oRb5olG6
w8lDD0w9az0Lei0dIJx2dXP6yn1kXRKNbQeW8wgwaDYMHXV7QbL26oejatAgTI64
HLu+RyLlChLELjLX6p6vj2xMiAp9GXGCEsuNfarxrTF7OQxE7UfaliMgl2GnjXrZ
YlPtlQZeUuySWX1K0hjiCWP50uuPWrho/qZCkpa27ZTEeyx+iS5D8OFdPw9dNAoG
QbBaA1HwHCBy95HRBq4VjEXCl5z8YaYJWoLTP6DbbiOXJz39iH61XVa5sUedVQ1G
xhoB7vvlLgU0Z0X5OgoH6LA4mRh0K7+MuCF7zYyubT37jKuwsUC/wnl2gUN/ns+m
qN1YJtcw+6ZPtHDt8ZQcKnxVns/EARen3HqoQjnDGOzC/5A+II7H9Q4W60WqQmyv
JcIu/FCKhg6X5yqj0EjYu5wa2IfDPHCYSLaCJiTwd4IhdiWO1c7V7PRwd84kiLlK
LJmG+++vRgLT6+cwyQuvMwTuRz9GBxB1GWaXKhlzCvTrkRoBDLpSkXk/hgkVzegt
9Vo8PJXcru+nobi5mtSMEEOpjr8KQGtyTglfrLAX5tceRcCBU2Bl3dza9/il+8uX
Z73ZdMFbQuiVzfxWshu3wtmjz2Tiwvrt9bmzGj//hgEfCGerPmtGdm2MZTN4I4ha
LL61k0aUu16ZUnCJdv97FtijMB2YopAVUf2XTZKKc/KYCd4M22NuaaMV/gBZ3fdO
yc11VJXBvh58FY6plBddywcY+0OOk2FPsl/P/mydbfLJ5lgWMmVUapyEMRNS3VAD
IkhbGnE5yW7axw7yTFvlctMicvhOF7Gc9+V8wVDB+eS0hv4uxYhMWQqQKB7QRBOK
jnxTgJ7Df3GcyrgNMgrK9b5peTIkzexE5sdMcdxgLOB2aRWYfuQRnwtBnzMqUC7j
mRVaoIutuWTP43FjBsSNcKB87HdwiBEwcCaAKAklTBx8MXnAcpAp5fFss1xBL/RK
knnY0UDT/DsNfT3ykU6KtWaKemZ33qt17KsE2xZrJHvtD/Za+kBqzwgEjiRCZsWS
ulbsMZmCcZ/+6beGIZd/N81eR+Kywd1HtCSBJqfQnpxggw4JUW57G75omVlwZPq7
gPAeiIaq1ceL3M5RNL8UcmylQjm6s6z/0SMmD5GsQzsiHlXgjKANuuE65xPYCo0z
2ALQDqzLmxV08UQZu/fKu5+ocF8WOc6iA40bV3Pq0aDm4lQzIqNLhqS4NST9L5EB
yV5twa1DotKWnyuqL8f0PCtPzGa7O/+l6Q7vKitJsuVnPpRqqHvFWk/NPHgFUQo6
7cdtj1JnfstcWIj5DWns2lHALQG0p9OKn93OfC/sw3GETKnRyghzcNaIkItbQurR
MCI1W9BW7Me6zQyiQT+taHOuEeWcNAiwsxZigTvwZ4OJD5jKmUO/U1emx6v6Ddka
7+hMcUDp9iA49GktU69ylPKS4SjfYEzXujp3s5qkWxY8WcS0PPaqt+tNhd+tCQaH
ZYzCnWI9fDg4PNevRWgwKgHm1RoHPiedWL5Jwv7176t5xVXkGso2B4v4KE7O8ScN
3GAfT56BEgg90ZqvSJw3egEP2O3+6NY9Xh5vYdkf8LXa4TPAOcNQct89YIjHHFbw
7sBmrq1Ghs4m7lMv04MHO5Hjr/BcYr0JZ5JmydnCAQFFsV4XorMK+JPwuk0gbvA2
8qhxH16xuCSeOZWrEkyb07OJ2OSoPWqzR82sBLNdrdjeKpo/sZX77G37wJOesiRv
96eIiv5wvxauv3CTOB0y3s7E0alby7zuTvTFXefrqpz58dBE3phxj+tBjMd+3zAB
ExxBt4YyDqEmIUAsI15yNJGYtMWHq7ty4zZPT6qF0qJpNd8XM6a1+ix+46ExrBMC
CsgT6GTixjUIxj47M0T81CQTks3IredhwStN2kOAtZ7P6blyV8xZAu9iRfkAmwwc
sJbOF08hxrziuseGWlxmHiPh6CvsrbSH9b7x5yQPmytZSXHsPWnL25tJuf/eYb3T
zvIoCgQcxOh8i3NrCPb7z02l46eg6CukmsbJi5/XUbSQW2ltfa0N1wF/dHqpxYZV
2QA2tJEi4SRadeYO1KSvGeq7MssVKFUdkisc36KbBQ6cMgdDR/6yZqrZYPBqVHhp
BfxAb6D/0ylsZFCRiiReFqJVXMfIdjxdHOPDW4jBn4dNUFSB8RyIy0qwRNIcOfe5
W+GK2bRb0pSsQagUfhAjJkPQuv9WvKcbz1DbsAIHtd/1os10HKl0CeXrNWR2YzsD
c8ATWeFcOVBEB6EnKXvEm/JK+HojpADtc4Ncr8roA/iJ9GoY/u0bGC7MPtgmGzeI
yZvT9cDsI1pLXhWbLXyw+S1IhmrDkKMPQS5rCRJEIjicXRli8ssrODdF+0tWJMme
4kr+4aKBv9xhux+H2YiPicI1RNQU/s2kPRvhOaFUgprlMD8foWuwR2uLmBXLrmWR
lawJZPuFSaeU7FVqtm1g01Qy2eEqkALyP2DuIkw2rgC8oEQGpFYtj8weowtmyRMc
1lvsJTyzjhSCHX2JivPkiGoDi1bYnVRJkvdZGMSUoTDoA8D1rsKY9QHx0WQeSiL3
fDHRjMrmFo949tM8UWhJmEF657IGLxfmSZ8tNWLdsSv/Os5fbrCugHHYzx50FrmZ
6yqATqNU7gRYQo09B+twdhJdzg9/J0fnrSstz65plOeeZde3sxJleo2/89TbOFWe
bhJSZEYuHUcg3lhfbroNgHzJG65XsLkKJ3teo2j6w4Hq+03aa75LUTWOzK+FEh1s
5Ikkxg1x369LIflV3STHHjwC67xgVdg1wXrcsADTyY/+HMMuu8XW8zVi/9fPUHmq
FBoaPKstoon7j/LsKQSOEe1/3ETxaXJnrNoVl3axkSbSNzgVJeMopxiybxIhUxt2
OLC+P8+FMQNsZPr6L/pRKoInzmfAfFhgQYrJEt5AqBN6Jhs28OCv2NlG+qockwqW
o2k352y3kuQN98ZzEtfL3rrRVw20cei4zfrsaxfeW8QE9EZsyRxltOfpB59k8YK2
GlvQ2yLq1QzMLZRoPKNn1BpdDGU8VK9SBllOx11Kv2bM7AbUFfiq9Qgb8Yf+gwUC
aCsj+DTfbP0Ox0cwJxVs4t3KYryl6yfNncjR0gDFZPrnZ7DuEJVxHxq3dCjTTdeT
SMkv6RHdm0g25m3Zy6teI01JJqGWFRixDVU1aRV6JAFtqzi2QLEXWfuL4CH/3p/2
D5jNAFl+0xfGY5CaUlVC/34F3NunnZdecMq1SGh4leCeRHz+jLCfmT4O9e11yFF+
/drM7mBJhacdpYN89ZCu77KwitnfFWY7+mRgMnoMADGsqbTXmIM6GxDr0u//z5ge
Ft1L/jyLAEZ4mfg8L+WvWSh0fWZ+haGHkPTcX6om6uZp2OXn1qPX6ERKa2gVQ8mM
vbat4kq4Qmfio+FsD1ry2ZeaGJqFRsCSV512yxEZ8iqKKEN5r+gnzkimhK4B98V4
oK1pSi1ecIYN7+QnVKqEOBDP7w72qteM56XZzoyS9atJOxmeRCj5//2Ci7ClqlLW
xpPRcyeSGhbpCsDWpRHp5VjG1G7ZCFGChRfM+ILtDZYn/WRhTk6ZwcUgzl90onH4
LC3O8CRpfJqH00B/zEAx37hvt3LAtwpt31gfPxrMu+SSuDLzOrng8xa9GELi327r
XDWzeyHptNUv26VkJjcgQFErdFhZirqx0779OkRcy6HiHP9qX5fhxCCoLAwm+Wkl
BX6iu0L+zP8sJxqtr7++YOeKSwO5KYXt3fVnsP3YwbUpjCcrlzfExBpAJU2Ee45z
o/a5K0OyrKEvr55036OtyLpcb0o0/mg6IxbtbycYarA0Tt9BU8olq47LLIWLDksL
zaLlk8QRbr1+eOICKi4i+C9JtxilE5nd9tL8xl2zqQZ/nW4lMxVt2s/f4Sh+w2bp
z6CZ8uoFSYG7VTCiSgfPKdd4Mqu2HTVOoCoP7POn9r1DfSA+ial/+8Dx4Qhpt8X5
Rt+O6m6ho8gWQG6Deg84cIB6EsCaXHNsarUBmu99H9CVKSDZPibFbPLttRlMCLqU
qy1rRV36akG4oVEIGTv8QaCzT/OMQHaxmDPapma5KXOXMnZrajVUWH/+1UNaRayg
AWpsW5yK1NB/6SkqX94GY6spCWKdLIabG5aHfHgygb1oH0nvEvOw1y9alLa8vIeE
ZgDJAB1ufzX2PpIB6W+TixGan3s34kzJainod/T1tn/ui2nqI6MZm0lU+GW14ekF
Xb2Qtv9Eu+FGeQNThcmoODl3dlgoBopzqzXkTvzq+7PDkuy7aMpCTYIWBlOauQ7P
mt+wzBblWeMiJyi6grT+Cc3yV3XbZBkNAjaQapyyloQvi/Im9777YLmaB411lmgS
2372oYLl8eB8C45CD+KGYx/Ndd8q3PhhpEJm4QeUn2u/s/YRGpz2FE7IawGl6Wc1
gJvOJEYdEZYDASbgRoNAe4nKMnPKkTx60jI+P+037bw7D/1BNQmA8rh4aywdWke7
Y8A2dhwi04dDMopLWpjyScAHx6T2wMmpnEtpBvJAlrhjbfnNjxUXpfohusR8Jbdw
c6hvaKmAGqPA15oFXqX4b0UXlne7lqiaChHPrZ00m1sL0T2xC3SqqTuye0NDAydm
bESSG/ZH+kVb+pNs5zBxXuWb8S9GT12cX4+xrOb+3QiAHPiBLiCuuXh/GFYRLrOb
AICjmQU0JjuFPfVw+7S56nzyjk5J4Q+wz9O0G1lCtWz+c3VhzNFTrMGPJHg9rW4T
9zqtzETlNEspgsdb4C3MrPltJ3y148go5cwv5rJkWfzuuS1r7wkCck41Kzwrob2J
tWU+jbi7TbyL+PwynQBVM6trRbT76SB3N9wX1e0sHU+lmLtibV9CQHRh1bV1qNtd
qQ+2pMPvdurdzp0eASVnzkp839g3wQ3RhxdMJ/SkOrw5Z+W/Bvfjda0jA5Vh1n1K
pW60sR+o7bDUNnfFGTeUk+6hCh+FoBJ7uTqgL4McXr1z0EOp9jAMhoks8u8d0YP2
PDuei/FJve3+dsdQ3gG1zjOp78Fw7so51IaS1/Z5E3DPSnWcdYmIsleTmtz1cn4S
lfPLlg4+lYtRBgIFoinV9eumU5UTaAeRxZK0aXApFKs0drHYpaP6hvkIDDtpo/U5
GA+xKoTZxVSS4dZIrLY/QIVPIBFI24goS7OcuvzSGQqoBerEVVaNDWxnvUdCpnNa
F4YOx/zwnAp2Pf2FLS5TRgchSqro9VFvHUFfET7LKOq3ETv54voYFa0n9hpGeW9D
zOrU0A+ZwEsK+m5PPjE6rEzXtxqV56wizetxt3jlUCgpz4jvyLmK1dFzyepWK9Ri
D+c3TtbugNe/Lbi35nKE0r6kDXCtW+51sCxmaPGGRCxzznCI99/51PswMSaS9UDr
ptvaU7/J9bYikscScds4m/FwSV20sngxze+kT4pqpMSgTZ9r3WqcO1WJXWh8hgqz
T/fnVg2hLr0YDNvs8pmmbcLNFlDVw+x8bDA4tec0opj+XuUBvB7qq2jS8FPYV81Q
7LL27CTeHT6p6Ltk3SYQqk7eh4Qpz1VCzJA8+EUE2ZbjHPE13ARddPcZTStqYI8v
+D0nBDU30DYveJimHKWPnE2MQneyQAc+cccZb64WczcW9KQF+qomN1lZTDSWY7fG
4r2WNmB+tHpBVSFMlyzSpYJ17+djb+jA9yfqclqGVfeEf2RUO/1drdxptej2YpNt
DdAfWzkQp3Py0aa06o4uPhksh/31D0Gvuti63eQYGab9UyvJlTrYeRC9d21VVKlQ
E/qd9RnlTgJhDcu6sNxVPlTLyctWuAHm9QWHDCm6oPz5D1w2KjGIjvVqOYrjKZFt
5Uj16MlJvQNLCv1kJmZIe3nMLsiPnI0g8i9HQq4iXepotcl07Nalrv/vrumZKgNV
ExSGpYnKj/Pvf3MTwH6z7g6SL1bUyvyIx8lYmTWaF9e6Uycj2QLLNbhfbmKx3CBx
SqGS2zK2zUpGXo9t65Y9bOJGSlSGc//BAvmIRj6c/excawDu0i/SW1c/Hp/Zb0ka
hYgUvmyQ1nK1pmQ+/x8N3XX9txmZC8KS43ugZiSZji2Chgf6Wq34v7WdPCqC/00S
ldLo3vyBfaz7UEtBwEsuf8Wyc1VFSufTooKdj28k3YqVCzn/PZAIIBY9lrQfCJSH
81u2HQP7RGCXp8lU4GqmAhxX40xKmQXsmZNFtEZRLBvCE6jiz7iZO6v8hjRb8bk2
bFHk/F9xVU3g+3xhbcIG3ZqZYiVqg/z8md65m7KltMOqoGCuHuT30tRCPpd8xuUB
TO72rwsUQH/6Rcggr8wciEfk4TCEMRab1aCo6ScpA3CBuIzi0FpCb/Nsgxp3Kpo3
cXWUYjEuLaJ07iabc5f8Qht4MW6wf8Nvi9Hdy6hQ0WJeAtjpIvdLd/TnmsDla/cT
x8p8C7mCIGMzsZs/iSvurz5wQYiucKooWi+Z66uGpjAveP4MIhBZKGtmJebVJltA
zNnDwA3NrYBVI0XM1OavJnV3E1BPIw/5fwWlcKoTPubfLaseVM+Fw6tg5i9WypSQ
8Oub2q64E9UZafOUmO9lWICSsqePk4Em+OE9b9cQUbBGnCCycw6RNb78MkX+6lff
x9ekG0s+Os9C3zF+m40Dt67RLpm8Y2hLOtrLjHuHhOkGD4wIW1Nz+Q5tdhOLFz4e
HbBR28Q8Xl1i4Qjm/acPgJ1hgCxQUa7UYpiqqzmgKTzcA0znPKm6s3FTZe+8zdjg
h+J21jzvuG/wJs55nRABrfJAc9bYXelyZSGUxPPW8341TKC2JooKjMHpr4gz3YHH
y04Oo6c3cC4V8LEfuBuDYiKttOdOEk/izcnQGQVn25wYZ0H4cUEHWQjFjtsIL7eS
zkYytDkqD4JJfgESirix3RZReX2xIn2ivfiQBX0PwVCNHYe18iQPKWdtrmwXIVS+
4tWWdYaIt549A7U9p+XC7RfyUCVRH4ylqx/X8weXl940zhynCle25r9TM1nMDiTu
22F6LqO4+5DZiRXUWdcUQeLcAoN6SxZXYHMm00KTHsIq/r6jl+yyId5ldhPpkFZ4
IdcYISRc2z2+l6aW58VvzgnXmhOa+tjk0RFHSdIDDXMTXjtFIWbmVHUb87KKbMiD
zce78MRTjJEjW02xh1/xtG9UivY021290ifLgr3eaUp4XGc2/JeZPQvyMQbLnRe4
FGmCRQ2T4VDHYJWi17RXAVp4B2sd9Z8wA/dzvtLQ0cp06eMfgVDCWkxQRmhxxZRc
dSVXk6Fcr3UukvZwJGpZAzSLImZQxjMorBVl2d7IWsM4KKBvc7MoLMWGjFgc+J3i
V30I5mjBRYvXgBlZBet47mPRgCScSdFIH3oLQ91SEG3LerJT8WCNywLcvQhytI/O
4aTw12INkJZcj5VZVf0xKQY+MUBZT47EjFb/frTPwr64TehAZ6fzhNM71F+OW8LE
JnKa1MzDv7J9gDRAqyyFB36aY1FmCdDLYnSabX4JBOdKgrVQygc1664KRtMbluPK
h4IkCCDjq5TE8m5HTi60IIA8JYgTPrURdoas5svAXY+jmOHzcdlQ7wO9OssFmFkj
UWv1ajYE7j2LM6fu1XaQ2exAhoszhPXoPwgF6b8Y52we5cRBm6qzR8cpsnfEJ9nm
sbDV49lyDRr2NJMhMtMFzfNvg9Ja2e1MUwE0zQ+zJoty6UvtCXr5NJz7fU0Z6uWG
RkRQ7YNNMxo0KFijT6hL3bJLafoQXP7FePBY58FGFNhcDKdEEN4irSwNMuY3Oubf
P1404hzCejH82f3XI8ZYi4drQBYsx5hBMzdU1YJJgkhHAb+ryBupBIDhwRKxr+1c
ZMWbS+aq8+HZKG968lSWrsBQGJwwQL1Ik0Yua4mqu/tQSzQ7ZwDTuHVntEe5d1c+
zr78W3i+1rIaMQ+af0af0rEY5uiKg2ReO+zarcPAtYfAlgGJxUflKyv+U/6teTfl
06AC003fABC6NuSQftmmSIbm6R359+TpIYyNIqdt/UHLWThX2MHQCgvNS/29phD3
G8d7CsYy5TqjqbqDWsH4aiBY0C2Qmq6QtzRpT0O0WpWwF3wrbOS8+iFo9QjbD2+V
WJ3O5KMlVQqoRsD3xIJdYxAMq00dCXyJu38UmCccYucApWyv40rJKna4jesWLuoU
2hcgc1Q+ZWjuL6i3arsFzQoE0/gUDKbYAjsDmYzdKkuL8BfmzEVeJwHrDH0Sxk73
8EY/TKL6XxOUoI87APYGAFv5YvxEAYOh93taOZKmI5FjPY6Xh/x4yuH7i5MOux4Y
VdZ/vg27hx/AxjB5BlVaLxsAbiH7moWEb0uHi7rgY8b+dfZkeKq6+0w5E38npxes
iKXF+2JKQAqEHPYEnBgdRjdJyAG5bYn0l6W/5fruXLEGku68X93cPifuMtQagfDq
vT/s/fCKhoOED9bFw5i8yf1E5J9tyoEjvRL8WGSGAkc/wSnkxhN3sqevH3qVMnwj
EM90mq6mx1u6nUTAeXKFDGmr8eKPYY8cQEVG7V1QOCsTh+K1uKMLCkRBl+bxjKvI
JpgWUmLs68S+MUIMOgqb8TbtegsUCi7x7DlDbZ5pYCg8+Gu3/WXS8TQcOQ+ZNR9f
xxZUmrulkilqaeh8mEEr4/iWx+TenWjqLBfg6aHdc5LJzBOE21MAOUS75s0gRSG3
MRVQBlwWps0g2XaCwqPYAwMiDnQMIPmXrJQgHHdiQb3/UHy2gwVwobNetti4ObA7
BhglKxcI7HKEglelJiH+P+nPI6gD6bBd1dY2zt/GkPzWWr/0oQMKpgnSzQg+8Tto
DKVxzpI+ZZsCFax4xxhDBl8Qswww/bXuxyxG3nQFCJgMK1EFrKB6n9nlNUfPM2Uy
xjWGPvKfX2HXIDn81NidRmSAGGrs492H69uQovvD2Foezx/sEAg7JnRIypXAyAHa
kl/SX6BvmK1lLO0u/pUEuiV6McAbcpUqKeqZ56rtRNWKCV/vJ3W8Da4bDy9TLWk+
8gq9MP6l6jV4tmjD45NzFa1yW72VJinvVj/WtR0UDAMSyktp082kuNxYyFehmETW
jdlZ8uGQ0/L4nj4gX5H3yRc5j3mklr8hiuizT2APx09NZtQCVOdbfSbnZH7R3+MH
0SeUgvfF2Je5C6u41G8lewpdiPDIRHzSyNiHZpl7dOadr40qirPRLjGg/8LPOgUf
mnJMkDqfP/TSvt5etG/aLeRngUa0cyC+dLCzLnr9Gee0FMAH5ZQq9Qil6XuIcGul
TSRe5FAwIIRovEbaLDFsJ3Q3R9S6IJ0JnCkmie0AykKlbdwy30Gi6YBUgb/YsFkb
VYgwIoIDIrTD0N0X2wWnnSIsp/tLfG+hIh40Sheq3ZMyRcVbRjnFrSIVpOsU3ytL
sj4rivooJf+I842iuEbTf/vh3rZYcpYlPNgaBvWyuhf06l16kt0cMFGqPZ6yiIfM
yWv0QS8Xe06ICSdc+J2HGSOMP6f3hHjRzg2/f6o5Loln4Jmrse2+LnuX66guXlsl
9BSRUwLo7xgMup2xpplKecJc2EjPBRQNsYucGSxxAi0/BwqZ0TsO/07HPp58Q1ZD
I5WPg3ad2uYdWJOtBCuVWsuUd8RbVkEicwuSzlxCzjEkd+Ooyhh8TfWwbIBCF0h5
bK5JSBurmNL6HzgyeUDIkZpWkDv1loNfwpDEBkPG+fPi3zQXHeLanxXkU/DKYum9
UKanXYK8mSSlsqtOtjAI7XUbUbmpFUkLfyHkaHSQLlgFZdIF2k91zYIgFEfVVTm6
gMnTh/Fxtfmej3NqDpDZfUI6Ouiq3r+eYM6UAbA4oeOArsE1vjDygVxYejfBTTRX
bG0tFv1wD+S4gznRCG2vFUDMsrBJsIJNqxUexhgT3weui7ZTwIbgLGLIWZT6M4b4
2bWpkiqcV1nvO+c4P8Dm5RGk8CdZDwIH1UAbqzTik6XleFNAbpHKqlatKF6NKUOk
jBN4BD4NrsARFXWAdSzo5oOghpJmfQQHsh5sJcjVmcOjDuQDzPpO96sP1UrqfzB6
2Y3WpqKRZzdx7HTzoK+wNDhNCFTZeLTyNb1gztcldVRr6UbgfKfEcOCqq2YuNsxA
210tosbhLAueqUOEypy8TOcqa2URBapxO5XkRSpW0tY9Nv3LriXl8ILsxS3PxCZR
9E/4afm0cN6yMiZa5D4z4zO9llSK0eX3uW7QMLKaQcCW9nnwSnrwz3+g6ht2v61l
d0gGJ8q2zU6aAZylWdei+ExQXEvld/27DEVTEYwsnN+jXx9hMWCyHuU2GJnXh3mV
lzpMsflSq1kh+vtrUNaACvdslBb2PTSHxL6td7YdicImExkuzj+rRMeUJvnyQiFH
OG4vJDt/5Q73tukhz/z8QvMH6Pwcf60iQQL3FCxnjzZTM2vRt0+4TaJ9NIgkWuq9
pBx6uH+ieWNZmcAoiba9mBsteUYo46tPclJjxQjZfcvDv+HHpcQPwxvjvpf61LzN
+lHSxT8RZ2gB4P0+LqaET37IeOI75oiCd7FYvv8wcXgINZr53OSJdGJm+Ungitmm
2mpnef789gXAJxbZYWPwxyQLqBzvw2YAaUixvHjUusJ5o2mzh62zvzU8Uf3ZjunA
bk5JtNBJiDHylgtDCSeGcvdbMmHHnHsRjV1h5SYTCUldSivwC5gC3aIK6wLq/okS
uC2fcm5C36nFRRVMwOQQIdeG9fsRPiCCN7kUt1WyTkBIOVdXrFl62WkhfWRHykh7
dA94rjT4awSTXdQ9fFKBIzZy5uWKZ8FIeCF2ZCgxOEW4X5Al8YJZwvcI//pbfaKZ
vzW9mfWnI7As4r9Lh8NIfXu48+qhEVA9xlFUA88YCfsFmHxeacmlAV5l1dgEaTAQ
ce+8RRTU3XYqbw1zBoAptaROFiyCidBdmOvd8MctAQ1FrPq5TK2Pr0PqO7POpbo0
XvYU6ysDQYTztAsWkgIiv95mvOjS8nK3sml40hnGNyljB26xKsZd1gC1JlNlIMXb
nanOooO4BMteeI3s6Y1MFpFpMc1sbYnYQwUy+OXI+rqFeeUkmmwnXfjF+JnPWVbs
432LqFJyqbWynTjRfDJNzpWZuxonIw/H+4lIMiSCuOxixRmiPkkASEzWpsfP0PnD
vjeGfbgzg1lA7fj/L+Mu5lCH1KFn568BhU14TeX2QmIXSRYstVZIqUo2rnkeRH78
tSq2KRh4f5o/V7UUJZzgo/EHHjvMUj1s+Tm0mD0z2Oj4MlMsfu/SnNNpf3C07AMz
noOiAOWXTSszwVBxN1427vSMDUJEl7PiWsMgOMaVEMtOOmQrWJQ985Ieu9nR4dTy
BUjeSGTTYV9gSFeZyUuNIWiqrsOCnpWauo3ix/pcvPwwnVDGMykb2ZI3s7YDPYzw
I1yXjFlPCQ9506FgN8Tg+kTThajJnanZq5xj/0vWIF47EhwgFdBE/+7drv5GMyoS
tZZkRGXUQfUllO+r2334hhTybq4gwI2aNQlZeYpmLub+JAa/z2TH9q5XEDy2VNbz
VKcgqgtlq1aCs6AaoP4wcFnMiZ272osRHkM2XMb/eqxKMKUpzMXnnVaiIUdSSKdK
pi9q8gXiuXTNcy8IOQUMm1k6RjJCkDWh1UU7lXL4rO/XyDX553GUgaVOh9XR5cSh
ff673bX19qCudsxD8aAIgiCje5Kd8QOsAIl6YS+duoqkNzrRit9cvHEFc4D4GGeY
0wgUht2xbRDHW8OeThwR0Su6Iep9UVPyAoo/6/93yPorJcrioUm5ZidUGg5MFWoI
AbVQeecaK75shOWpvG9mU8bZ7TG/TORga2iahaoOHzDI6eFz8KDW9uCI6m7BkO8n
C105wkksDeAN6NC/Ll+922jpZNAV5rjnrm4lME1vhXAp7dyXq+0mh77rKovtMoH7
rGFi3fDkw6QwOzyocqjCQHaXENv/3/3gwxGbUYnqQbnu61Gw1wcZhjE55U3K9nmP
u0qapUKJ7rc1FpK2SNIk2j9NA4L6w+9+Jit2Ebv9BBaznx7BHPWuVhw3RpTSWbKR
ZxA2v5ybAtyEA6zE3hwKtDXyDpskjjXxoU95OlAFwr90K17OvJB6C/MUTppXgSRO
2ogEH2tMv1nxkK4HVuEql12nNYcx3+zoS9JFW3x8FB+kwPP5B+PRoT8jyhyMiJC2
d2KWNbR74mEYtqjYq2WK6Y3O8u5aByYw+r08lkY5r6L5tAdHJu7O8J6sAXQoAGQv
MMqQ6WmoSzoBbS0Nw7NyYAGdWswxfwEDYi+zj1m8LqyG+P4uni5fUJy/iLGpkdiz
madu8ojn4JNYhpz9jEgm7jkISo0Dpdl3zWRVIzSx7ypSRC9uBzaJZ7MElwZYRe0X
CS3BXMChBF8in2C6Y1Uo7M6ZgKx5c3zw4c2fKEtxiZ26i0cpwXjdzwMJB5xDMwhe
zW84WQ61BBc0Q9mYRHfRYiOzyu9+5+KlnU7LaqiIRbeVWFa0wPqmCG8PmvoD26N2
Msqg/fU7TyVOTbP1+D/45Cv15L+5Toh+f2vsGyFSgqEHLfLlLJNALuc90yw+KN0u
MBhy+RqeCqMzO3c3MLypSB6c09RWgKkvxK8uyA6PDuBZYXhmdt4WmEAhgCT82ciC
ebgNumFM7EpWMfPbj2joMJ/8un+AB6+rcibD+hC3DQQVH6IiR1HFNMQKm9j62PPs
CF0c028Iu4KNtFnXnLT3Vsilg7+XMkI3WZuRpnU/QSEt+bOxu+re4AMWa+hBdiwL
jpFc1dXgwrf0pSpQvLnobPUzhmpJznn5u4UnxXhSmwVL1e2yVeJRJ+52zkVTHslB
ulGEPFWritM7ytGqxhl6qh5pS2ITa/xC1gjcufRnBsOIvRyt6Gj4NlQ/vmo2okL7
EDd34HlOMQ6Ttdb4dEkvZUoQDGus99z+UjEGMWrMheDhdmTsvKFMx7zfpuACqk4X
UtFVbPCUTqBN/tzopkLr+zXJEcNp0FbfzpabZibuipiQhGM0gMa1T3Y76A1JsgMM
qo7IaxeyS/bmf1mGakVUB2kL77oysN9gy1I+bky64pja4W5rZe4I5+s9GAJs2Mqd
zt6dPvf0+Q/fxu7CwxRQvsEXyorKagwxKS9R5YhOhRUddG+voWPMBFkQi1QHV21W
u+GT6Y3AptXYHNhNHzVT14em9scJXifwoqSdhZaENXapLX5U5TT3wgI53STvUlOq
pd32C+Wd9zykdcWbHcWPaaE0ylvX+KV+TU4TwDTvyHhRSmI+AiEgQof8VPBjKWe1
CmhLXj4sfpPlIjSiXdOvbtEX1+aBdWzvZGQ24aboe6Rgbe0e0/qZY69p/TrHRMYU
jQbGQVVUwVlN2KVN/CV1R/xZU6UllDYR9txjBYHkg2cYkfZQ5b21E4oF6c7qRMFc
TKmwUQUegIsMfLMmZFJqAzCCRnIgmgQos8u4R/7gAecSnkbm/YIk5HL4ciLEC3ey
u38yTdaAIR94SYY1qjGO3B/dYAHsgAuIBaw3plsjtbN7dO+ZhtAvUZfelVhLNy1G
FZSMFHsUjIr276aIvvBjFrSuWG4N/yKXVgwA16LQa4QiB1tJf9NIo0iMMYPOuVTO
xqSGoaofrpbA8IqTT32uSBbaxrijBRxicouNVxILxZb6o4PaMvXUQ4qqZ6v01VI2
Q4gzY0LVanWDW29M4EPUWAZxecGbrzelY3hAWQFD0dimi8szZa5mxEIAwR/rbOXv
udBTJSUcT3QOXNFYVJ9KM9G5Mc/aWZzvvVJYa4xSmHXIxPtRb2rbhJzMncLV//4X
Dpgi59D+3XYa0OfGqMaRnb8Io01JsLk8MRwyfzLOFrBt9nhLBoeANgB7SCZ+/yO9
lmp7mOG+JI/Oo4/QrCLAPRTEyE2HLHtUxHHVnEglPjmUJ2XFzRGT3XZrtcTq6Sx4
hxKqwz2+ibEHYOMZnUOf4u8Dun9IgfP6Q4Q9vHwP59DQwGrv7rZFXLuOPxc1+yJb
rLx6gwJPW7wv6UR17m2kHBHIev9EESxgzo1QZQo70GF82E2D23zUqgk7o96Uegb5
0d2L0HwDFBBXR8kN6bhRc3SnqhP0MGE84wenVn79+bPzIr1K2/19PZYurKLuNFT3
kC6qxqLuOgkTBsIMjGaxEWv866LISh8bg0XOUH+zsOm4UN8sT1GGVEX/yHuO6BVd
pkRvpFxQUL5IreKYVsgAO1F04SqPdJ4zE7Q+OyAhM4Ko4356Np9b2F+JrYwZrRvx
mkfx7AO9hwQiDgnb8L3hEj/MgMaLtnRnZwgQdfZiCbLXTZrNdAYUz2tahd5P9XUn
K6gby1k9jcYmI6am8EdpE679/Lqm1yI+4/E9AEDWHJEeOL0FRtaCAbzSMJQHbX2b
NgmztvCl10j5TtcMSV17Wjx+M5cYEeFB9g4+eOUiye0ieYMBzbH4eGClWUZxUPDv
SwW1zJmmrFT4PNaEfv7h3IOtvCJfxG3ynrE14ke40gAma7Bom7fN9r7WRh8PTXqM
Z1HZv3Jd7pcgoF3ih76fti3QkOafx3G3lGSohPkLVsxPX1NVxVPKWN2SkrGIrokO
aBs2tNPRkUUHKWx6Arny+kSS9uOqdx4EzFYXsjyKK3IAWtfOFG7+zCqydNtVlTWX
85JOTIrKOIdCkA3Srb3bzrQACOeAR//AB7WjgX5cKDxzeEDYgB2L/TE7m9ecxTMw
uBz8css/bmNb9J0HRUr80qfqeEDGYcePVjLUJFo4cObzdqc8XsvxsdfBqeBAFaxx
9mkFzVdpH7Q3wwJstjos9hzlfBEGP3RQxeT7y8FVdbcxHjwZsNrMJav2eK4X9uqR
/Bq1CjP/DiAyIJEpHor+W9vqDGAYfyfvoNbroPp08oInFghcuOzEXnMhUHNVKk4H
Lpz+23r53dKdFOgG3KA9EFRmCifwn2m0wkkRDZc/oXgFyvdCMhKw3dFF2Oy/uv8d
fOr5nNuhiHVE5A+kwqiWIAvTkfk787O331huAGlwN+0RkQIq4CpZMmTWcAZi4Amj
Nqy+bQ+R/Q6/TlXmgnw4k4iYIfYxtBWYSP0YwjhI1eRXmd6bYTZJmt8EK91nQZJw
aSEIwjSYYZ6OndOcBZb92NAUYI53cJqGnfaZrlZBDZsos/EBlMVh1tlXljckmJqw
qu8G7LVzRSseefgYCR864cqts4/AvK+SUxHw0hrewrmh5zrVQXHErQiKgKiLr6cy
SyDIG1Hk3DK3ECsp2RFYoPLxOpe0OgSt4+KvU3VuSATpCEc7WWHaYbEebyLoIMq+
MR92VQXhtdQ+/aiP/ZK/z9CgMypc1KAfP2SViX0fj3J4DNTo5qwJvThraMozWd7O
e7ytu5odm+7AT7ZLF8C4Bx3V5vbBK+9tHMEBkcQknODYt1BRLezst0Top2g7Qoy7
pLWeset/KXpAsZ3z6azXkgG394dj9/5Clliifu51B11PjOjMiZegR6A12EvcMYvm
JiePEDRdzxd0hmJ7zfT2jyy1mIHAaM2iu7pXNKCdOB8b1i7/vs+jLesN2t8UKVwe
f/iKrX7Cyd3mNNIZtbU50Z9z+NSSKgIIRzQ9CUUPqqbUVjrgIrZB9VHjjANDbdKL
Ft0sM+ORX+whBj0TvQRNu1Djnd7+BQEXbrhXNFqAWSfk+BsK4EqWouJKi4BXb8q1
Jbp6+82bnxUjW/23Vpa/CPn/ijaNEW43fs8fy5TkJdRKkiv5ciYSnL6u0QbFvrKR
3wXHBTbUC4IUunsiV677WC69S1K5o7AllHXfH/yUI9WzK7MOihlcEe/NMCu2AtzC
VlRizL3clkGdJpjEy02NkfDbSEzxxp1S8p5zDGP8xHjMZRSmQBssVeBXzh6aZeoR
xt7UfafmGgkyOpZRlq4vpRN55EymwyuQy56O+xN0AUriMS+ZQlf4n2Qo5rhGj8mU
kjyrhOBqkNZyKHQsh6uPjuzmExeji955gS/it7d6Ddw+gLjS+ceJiuZE3gpXq1FM
lcj2+oTRWn0ApOGPztxLG9i5JsDBiXEBz8myv63vlkNFXxMW2ROw/80iduVAu7PV
KBxxCDWCJe37sIZzU0o+Ykq+eaHUJ/TNTy3ZU+BjWSTT+NMX3x+X6QQ9Epo0RlfS
BFEMMZTwzin9o/sT9sAuAvC4Hk9nLTI20wXQuYP7mAW/TFe7S2d3vHWmysMrokQH
K9dd1ygS7w3cZ5uh54sshGZJTavFMaA/5h3v/buba/6EarH6BuZQb98AAj93Zgog
CD64d+MKgddfEZIDMSzLVtpwYbiKQCyYKRgK763iYkzkky1DB8L/+HEsQAhRt/oa
pNCBQcpZbPcRuYJf+LDeKuuZ+WM49y/UbDf3x4ShIFwNfO98xEv5l+HJDLK/N38o
AYcet1rb4OD3cXkJfsUlb2DbUP49noPDIo248S/Jq5+qX5rt/s7K91qdMTnCdZt8
z5d7L9Y3wfMeMNQnPSAdcobGuk2rfdo8WO4WZQv84Jhu/f2SJaIDrpMShXWW67aW
Izx4cT3OkWhV3Ljyc2kqWqtEAottA9C6D3ZIuR2Agj5bt2Ik1hPjLdBh1wZmb7qj
pRtl5SkC5PSxs0A80rIIjTjPNVZt0o8YSO7NvtfbbYrjZZZmCGAYwOmP8wO4m9pf
T3EIC9eP7VWgIF+HuH1MSd3LVmeJo8F5LAaIapx2PhnRN8VrlAkFjzgzeeXnNFs1
l3XO3jQFZjwNSTHlVBUZag0yKFMrJi4ZVVN/zLCYs4c/HE/dBzUyQUUy7OwlnfVZ
yD1SSUHLzDp/v2WFVdF/YXzOWXiICXXVoLVOJWzelItaPlmSK77OpfXJjE9xaRsU
uiHnqGoh9haZ1gYEAqu2KP3lK3M6vomJdgezfLTygZgq2treaFj90Ex1NOYaZFhv
RW1F1ILVLr3m5ZZrGcl7+bgIuuwaSE1Ukva+LA1z2CF79qGjwHUAqQej92uLfnBU
IDAb2Y7rDMwN9bU0XqCRn8qK+f5eiAxTWsVcIqMvzvNPk0HxKmgsjCN60yOheP1s
WrNwQ2deB7HcJpsC1ba5woppr2kV5A8vZo2CHonbPUnid8hZv3aZRsadgvJe2/5A
kxXllV0hHJ1vmPXlMSR7pBJws6EQ/QOoflyYi6sXR6+7Oj1EnhbZ0+YC4b6PR60D
o+EE9H2cFX0ZFRNSrgOYWmMfqtgiukVeWZ+a8mn3g7IK9w3OZJ7orNV3m9q3jMCe
mYLAqqm/pXFBpUvA2voONkvRHNMafqxoVj/1w3MqMNC6ANTZh552lGhIvS3EjEJJ
0KNael1gvnzp1bG0eAFL4qL2fmNrVtdSvf4Zp49SpftJy8zesMpKOBJSZ8A9u/Ra
AzhEz5R/jn2Zidopp0hXbkLBKFJVLwW3/r/K6t6lRlG4CcWMfld2qVWRRB4CkE2B
68DLrtX8j94Ykblw161VPvQbdGl+YXgE3Vu7+8cT1dXlU8pnyxA1qgVTcBrROICe
QoTYCmgdywkNqMnLBx4+YThz5ulJyTXfpU3S3q7hpWl/0L82TshIdv2Eu2puLXD4
SyD5gl3RhZB244SjL/uqNfAlgMni4Is0OPBBreN+JMLx8HsoyhBqeoUMgOubyiye
pmBiVxcC+NhQzZSChrTnd/8hXKwXVPkBRsRKW049N35N91RJPJddnl0Bx1kHrqXP
O0yMrGFh42D8SsDzMjyXaTSzZRjSbHYCwIU1+Ym3dc7Pb6xY3sArepgKjRyAFYGo
yAuBAiKYYBe19lg9b/cZ23483XHhyBYiybH/FYaxUAV41qq+1OSij2htDg0nPuYV
QHiGS1PExOGHd/OF2GAcoxA9hbf/Nwka3Rtmjq6qqkmclxo9VCLxAEgMxhKn2cZs
rKLP8dmcfMLtwgV7eBAmxNup3t4HJnTX158Cuzfwxrjg8qOqLlZcGvAhXsEJIRQg
zdQfKPi7rMbdvmGouHjrIP5TSycVf6uNl9L5L41QzlrCRrvCPpRPROfWg8v7OFX/
Hx+KJZh69UdgYpWtfNFnVHJq+viLLm1oRpQaFUt6Ssdyn/aj0rIPJfC/vNeBIs2t
c4Blk0/i5FogO1E7yM6LUMoPzQFg/erVw2r1VwjIKVa0MeFM1jxeVw4BUGr6tDf8
ENlwrrHq8xzV1272ufwH3CJxf3fA5qxe+CgxamTEtswy6J21l8vJbzdJRLEyuejd
1IHo5EHx9jVhT/A3zRpmjFkAZRtDTefjagykrhQCmie2GcJhK+0dcTQRMTuxyH+Z
KehATnOCFLywCoSgk3Ck9Yf1WKH3ggWUtbd/YSOfzSzh24WOFwdsIwg4ss4a+WHk
mMVWi392Czxf81y2lJxKvxLhJtXXZge/Ca4Tfi7Iv5nWpWHEJIPbNKeQ01Z7J+S3
v/tib2C2dwdxcm/bYfHNupyyThiJNGp+UUfbXWcxSMTQhjH56WXMUoQVZGn/sPWB
DOpJeowApLkS3VuL9J6jokxBAQk/6tbKNE0DkVOofUqRhOxv60e9sNKDQ6uILhHp
7ej4ikrlIb4FrKJTq5jUr6G0gCimDRVV/7iVPRkrjL6Yoj1Unw94hZbUSdewNxXh
8JCYFlBmLTqDR5z5ddGibDrqFPHq8HMOjNtPXP4FCeiEpUBbr1SVd68Hx3mOL7xQ
sej70i75y5P4pMy8zxp3Vv3Q78id7t/TXJH140JDTwPE7eLWxLttiRvvuuJn1NDR
e6kZ4kzktWD/iQo2yDj0jbOjVf+rK8XFcvLUhgtXPK6UQjFa1FXEJtwN7xy68FxQ
dm6V0/h/IP13PidHomLE/xgPOdwZtxSROCWGLypkNYbY5rF4AOjv6B94GDpgpayj
ik3Aj5FGl6ubl/sIYr0jAFXhbupaZFlysJ7hEEnkyS3n830gsGct6bVEJ/u8WpBL
NrmKlKxJOLTwpKMSRmdfgbMNEgu3ghZUTV1VjZjqUZHWho0OeL6jyHtOsn3V5/lv
1I0bpnzUjnSMBjXkVsS1/DefOOvrb80MlvrS65hKiQabJrQiSUcad/EH4xfsX+8c
rZuZODsqCcjQPfFJd9075YfDmVYpy17FiBo2GvENJYooKrAMZtToxwxBRr31FuQs
3/LzF6DOok+PC6bQLrbut94OBmwsO92lHgXXhDLi0k8SaMpykXxkonj1wNOESL7L
1x+GeeJLFn2BvtvYna6r5VRU2tsB/yYjP7ABDlHFR9+YFyquFD/cxOgVCxsDLekB
RbtlBnh09q645aKSsgbqKu3wGxHS6P/adEHkrf43Ce0NDXksEO1Hcj2BIVjwzmNn
apnWCFOefT8aaZ3dJ+vdU/FBaNCXxtbpzrJjVHvAOvunYeLbtpZukEVYwyir6RoP
x5kjv5VwDsXIYo80Gloc+VIPQ0oBvPH4yZ021u79mOdAkVj4Q5QK6sNieli5amkh
5qT4np+JGulcfcNtOaLfgaTarjJ1Jga05Xi3keOkTDOqWkKi2x4cYUYPgaM2cWTB
2WdCyzJMuyvXXEk6JdyXDM5sVnFaTacGwAToiJSVwJcq/sV2HJruh2JyxU7iBsKE
39MSgDBMf+skqLiGyr1hNHwXhGO4+vsTW7L+a5tKF0vcpEdRLnUfT8F9KX7bwPGW
CCTKD38ZcvCLkbJO0qkub015Fc923Jy8/1bqNrUn6A7Q9hAP6MCQOFD17WSbyFZv
VIlZIoruTPDKTHzyCt1N+CsV62ogEhyC584NInxqHkFGlzhhwS8fL023gM+fqx2s
ZF3zCJJBlQvaU0ZhYJ3oiz1onOq8zwo91WLb0t/UH24fSjyAb6hZcgJtGMF0ssM6
SK6WL1nIN82ltyGljIwgJNn/4z5ZynoDaez/Ujz2iTedKN/3tnHofAWcEYvBQzpK
ZVeHMFnLJeCOu0LOSjyP1i0gOwO3ueZEXwL25ARTtEnboJdLltmcypPshNn5GwGt
QQKXXO//HssY/wWRzpWr4u2yIB41iJKxzQvItGLa6R+O3Uaoz/QVWVPGsuV3TMIl
irQ4RVpB3EWW0FVVRg5ufOD/nykTD605m/RzCKz5RdpGlzdv8oA/vq6phBBB92w9
tbTKkzh1kZvAbx8wTIaIlY6iuRY+6PTpmEid3BDPjc+RCPQe1pxE6ZFyrGwhDTcB
AvgpP7CNCiqBc24JGiaFVsKtI2ugQ306PWADpuBiOu+QkhBNyoXaTOrKqUP95F6c
6Mw8VywRA8woWWVJxS1JnHBSL5loLHSZnoolX49/bRtbZHTaDrkqPFgXPoQb0M7m
FkAAd8Q1iPzxZGOW4MwLl0SQgUSvRGH43Jz0Y8B9APY3vFp6moYD0hNd6tCchQaq
FwCMav9muJubtYiOYhSHwKtIWuNoltgyzf13Nei0SToub0V9F2S5i7R23g2XS6u4
/ziKbhN9siiWtqVeuKQ2mJC3UtE6k2kgWrcaQODFdocI8h+bbCBPqPhzqhhHDwzB
JEnQcVVfoIEWXlqlT1QOYfoQyNcUCF6PTp/WJ3fB4cKykuOuKMacmd5CYR2FYric
Z19bRnLy9JlJFfsktZP/ail0Q7DKg0dB94EO1ID/NVYRbOO/0gXY4ZywckaTfxPU
BwFngc+95SK2CiFnR9/0xx/9QuBv3lWZAD4OIDuqBAV7vgK9XyW9sGSBsoI48h3T
8c0F8uBCqYiCXCoFcBfjRoB+S1oXIbHld+clLBV7+t2foCn5NOaVbUDFFpdvUeN3
V7e6uqilUCn3op20+GIo6VS9xQbMa1KKRN1RV11rqxnV285enBglRuv/i3sG2Yx4
cwguvOeK3UnLH8IAUEZMlm0jN4BFRGaayhTtZgycsUtz3ya6TAoMDQG9aO563vIo
8kEHBAH1j/0A8uK/rsEbZXWm7Z4jkex7lOVShhOc4Xd/sKHdQC6M6a0CvXRYgtbq
UgJn7WDJub0OHfugfbj/EbcysaBfkrnmSSIIDvKimrzBeXdElznfaIhZR6GbN2WB
ea6b0KXnHM2U7qN/WV7X5tuawWIpsLjVwItlxxr+5BrbaTNbh2lmXKjQPb3PYqMq
eONWWOMa0UObOu1jaeA1ZaX47WgF4XNUUJK7cmM1UZK4KgFG1S0j0zDG5OsCgzv+
H1MEyowdnf2e7HB5SMv+HXPYNIrSn7uRu+RMdNpHDX8NocLsGvOchTvWawepB62a
fIrx8iRaCYWpnjsEfbA8SYg0e+gUYVw/XhubdfYT8Y+M5Y+IyqKv9chrqviuf0uL
IpS3BaMGDYoNbCV6VW8pdB/AigKuFOq5XQX4Bs0oqLi+IRW8Hw+tMM5kU7CvwgaK
QotDgkFoSLZqxSMAXqO4VbvmmoAHcgE7vK2qbXgD+tZJpOAPS9J132LZQsKKMvTg
A9Jc2/LFQBHzUcSfnu3NzgsT2S6gaNi481askJmq13yhteKe9q7ON1Cck4tv0jEX
Wjj54x1npbOPSWc9IfVh++nvoZvsZolGGS/4IqbJo5Nyb6fkwDaHtyZidss+oWL7
HRuCW7k2VDvBJsigvGJE7NpjJGO5oudD7UrnSRI6l7FIsvxRNSTRLk0p0HTGbq3d
mDbILXzDhx/SPidFjelvDzxAgr9ENVSjVwNIaDvkNpznlxwQdTe19L+YiEom69Yv
cACAZ0mKNkgJljt+WgRizlF0EfmHUsScUED4KVRq64oJl4hbBBZW9eYotofhskOH
sqPIPtPdZViLCmfQYpjnSmXMf/skrd6h32eh38U42ocbDIpYlnVtLtU2sU/Q2TFx
B8Qj6qjppNbdArrqVz5AjhsW4Jnh7rM9tk1uP4apobSLeLwRRESxdTTmxpbokJcx
/4XeLwr1Q3wSv0pvyixsoHQ5oDFIJNRZa92GD0UBsx40PJI6gRUY9VFOvPv3JjiR
TWEQakU/yH3xbZUTsC4uHNSVOewGdjOSYx2AlJ4ZHHo3fVB47CsKaMnR6Mc/tAM2
eAs32BoqEFvRFNMzT0UZzgwGEDPnmH5iE0kbJlr7/DVJr8QIEZyB/BWJ6PGQ49rg
X9pcVCuxsr3HQJpeDaraOiJIVxzOAACVgVgbNHUSn1J4gSYNyC+6cnYGwhNPXZye
7SW0qgL4XzTcJgWod5UIab3+MZUnj5oEFhoi1ygO8ChVRusEvoW2FCfsEbPlLzeu
Kl4Y5bnp6/gS7O5TAsDpFcl4sVnovbMzrsVyqnPOGBFcu8YWZgeLbHfgfiz1Ssi8
2D2Lz3vmzmaQO43RhuLSbJ4f7aaLGPh/psjyTGS/aLoq/MB6VtOFW7A022iW+r3W
dwpUQax5LUIJ+b/7VU/gaIpeIN8o4mRa6rxeCEHBB+laua5I/rXcY7W/mRM+HJAH
C3u7ZJm8lx9bVbNN62p6n8VfUjsCbq3/hTOZhFyDaX306QHuh9rqtC3vYdolWXL6
x+FZ1rOskycajNl2NiqociVcjqVmZZRhB2lUeT6VRajn0W4sHypKpEAbZkZI9DMh
RjREyacYvL+CXNS0gMK3+VQ7kVkwxSI64MYkGTfHIxDVgo3T1/8f+qaK5WWMw1xz
i6/VUINSW8Ob4HD9d2ElvXdCSH/rfGcOCmLYEKjcdzj1sInZqLmHEhUl9kcjEXtn
y8X3ALf2ZS7qNlcz2GMIWMvZko2/1NDCT/wtBmqIIe0+3ZlnAjr6V/ziZoN/PDtE
WFDGKhOxwr4pc0rbeY4U8+kiVxgFdC+Au8z32+GGwtYEZ/OtIq6LqmEHOw3POHi0
d1LdxiGELrh7IGrQBGIufGvFOdknUu4GKO6SFL6v8xf0LJ6m9M4JNTYA+coWbhVF
UvR4fdVaPlAvxXZDBIfMaHImA/tj9hQc7y5xxnkkKp/TtZkOKWd2FgBuVUJ7NKdl
jfHwexNQjjma9HMwuohK1nth3Z75U+C3f7Ozfu0UvwV28dykmmidwlklTlu3lDo5
tVvW2A++Sd0Kgrx29pUHMr1qbEMWcQsjpBhHCYxlFOGinfH8W0pp1mEx97fRwsDP
ID+MExP5cwswAzINCxF6ophaKWZuQGzRIxY0zwy1auNvMgM0nY/w+W7c175P7Les
68BHqnunWVANgMGPugNsjoP2OdEPDy2/lUUW9uD25RshlgeLGVq6R7eYnpilTTxZ
eFpNZUZgYuXfwOf8IXjPmR3m3ej06IAeCJ3NFa7J50soOXpWgFopWHiJfoLnshP9
wY335PfWjv0TzXvh9AkXZI/tnL3uY4Wjh2cogs56bnY+DlEjCsLNsPYruhlpq4uw
9jOEb7CSrEA5P++rug7y+4/RNl/UYDBz9Cf1w2JQE12IdpdVjD6HEkwhewCuncN7
+oCrOiaiWLAExsH8N2yV0nXdQL6ZU2Ja/dYmbHZIxMqJtLtLwudsS9yziX2YOj8K
enidMAHZLxSRFk8jjMujWduW9Pc8T6PKuHXEflgVEeka/UYpQWAHOY6ABNNO6GKT
FRfn2gqt+gfqU6Op+x1xj5CN4Pfve71R+xuhTJBmLlvLYlNZUwYj5Zr6x1+KHafw
hM7KejbZSowjLZWgUjktiy4px/Zi/sMO7wcr22iK7pLtT98zeCAdQNWhvn9X1eOi
aRxm7nHCxRZN3tLuVz+6kYWbM6/J6Xzw4OqBPT+cn1to4ZKc89b9LUKqPMOXkmuC
Ih2PmuJKpPrurGanlJSFr+RpzWu4KqBuz3lqEQg+S8ro3u1+/Y9V09DDmbf2+Way
0iWqnEw2tFMMLrZY9kGQkeUN/xE6wqoVAX3I9d8rStjUoC94cyvBX+oKrVuT2aXg
Fgg9i5vOdXuVi/Zd2/AKu63CZBp0l/iBZaGrHIJ8+eN8wSagpiuZvmUKBxkohEZU
B6RFpWSrSBjrH+bdady61+xtiLXZTejCv/j/E6YZHoRBqq48V8nr9fHvwcHVtV8w
47gvxa0x2DZzFdYsxLpgE/v/Dx3LOz+x8/1TbbP8MSHdxOOcU+tD+xlRNYoT4U8o
cSSUZpNYDvLcnbWCMk1Lwc/p87Vl56BpWIbOKITTzkOoV/2cFRPkgMAi1EIwFurG
Jp7zjGAjCrg349+Zmx1wyfgF9vkv/ZOD/taySc8vHkgfnqV/Usi4AolFhfdo0MHS
nx66cGq6b4li/LQuXCWqgBA0FR7LdzgyY9/tH2fTCr5YHZ/zyZiXun93kLuf/qvw
xa5R11mHPVtlWMiENONPx4DxrokE6zLNKAgt2o/g2sy2JnJW+MpEXslbaZNA4FJ6
bp5iJMruVOwUY5IQSZIcpEVhg002kBqm1kwYcFsOIVfQR00IfF2VrIhnDlpHOwe9
D7zLpvpcs7t8Hua1pZGoC4Nh6a5id8fpRjnj2XLezo0nDds4HgV3ucil8gOXeyQd
TdVrWi4KpzrpgDT8Pww8tTbKKFLRFF7LyzUw/HtbAffmCjqK62VGYhaIGYA8+vUr
nhIPA0E9CHb3UZHm6ykji39T4kJSvO/KNBUHCPfQmeoMzIjcAFfDmDxUdnFJ2zDN
kafYUicfFDlH27bcnS3MDgEpN1Z2cbnC+K1wN6ROXTBVxKQf9LWL2fKLdcUHDH1z
DifMEnZttYCyjs6S49Lfj0xnzgESyqNfA6uOc8zAJ7f2WzoHnUbTLlJS9goaYPrN
amSA2nfD0kHBvJdXqbb+TDw3gboAF8mZ38tgJ9G5tduwrTWJa8Am00WjvCIsauNZ
XPppdIC4rSrWJd0u781yi89oeCmndY9ne3p0HTgyroqvgrRvDzZRtXw0RkxYV9tW
pGNmdA2zeL7zJ8imdqbZK7/E6wB2YMnQGZcNLCO5rvknZDfAzyonYZ2nnxANj2PX
wDFrrqDwEcREJpi1QigHoT6RKsNlXbeFaboxoq11pgpd7Evju6K52pdryFkNumX4
19E8MccmjoBalNvM8AICybGp5mWWUVnWMNT+WM9F2d8xgBRnshmeJqTn0crnl+Qg
YTdhonIHTH8dUs7eBKVTUCz0/hfHrgmWjhjYjOHuXXR4VZiB9+DAJqBYz7pG5Cb4
ZtBOJzq/RvkYInu1InYrErpfmpdm8Ui9lArAjdfFlygp5mU7kGluS23aKc3efpvw
1zb7TkIOzibf7i8vtNi45tGJJ5uKDyozFqXjoH8+S/p9qT5l2NsD5MjZzW7KzOdW
DVF4K5acN9/ntMiu0p8k7K1aurqkTcO3DSUBGbcktefq0jDVbTGfn/oB7p2aTlWY
qS3ZpAwmz9DKGeRQYKhGBuUmtIqd3UCUoIp8uLPEZiLSmPPMZjG2GpqWf2iPz1fd
ZFONZSZ8eX8ZKcHhBhsoKUU9TQVvooE1BNZtPBJT53Ms0lkKHimxtv+y6WfoF8hf
K891MaaNInqYhpvKtx3M8+oTdeohD5gbHCgvJQDKVt0QJm3M3ELwBPAzgSYh1zuP
+4DpjFK5KolnbMgkKz4LpD5ZomPEj6VjbYhJf8/6QFgHTC0B2hy6M05hZX9/b747
iNl73LQorqE675R0799Jk2DADUd/RWsic8FQmxGeqHC0Gn3nRLbu8iWcUeQexnru
Nd1eyHWmUAM4kbz8vYHVM6NxMrAAyRdxzrBzpD00Ltgvf0eoqohbB/0qjEouk3xW
SCQKDu6p52bBvvyxdAJCBxKOzPS6ELL6PNoEE4eX0nfPK3P75iRoE02vLAhmWWwh
QOD6OfAKVfIjFCsTJdDXWyzPMw3qbmsB0svBKBCjl1W2nJeH8VHIMEI2ePx4o+DN
FM+uyQxF1sEmv5RNm4xK3e1JXY/OvGvRY34WZ/zUOxde1o50WDksjkmhc1k05csy
yjRYQLlwdGgDA4zLDsz1BOan+oJ5jOE2SLw61FRGjN87G1IPCM9k8UNoY2EUFRxl
qfNY5BB0BDdKw4xB8uf/O0I8VbG6nZmyKb9AZG4XiHHwYpWhw/E8vsXgBvX+90R2
UtD4mLXtapieUF/Vpgr4ybaZC6UPcH8WtpkBwdSuLaQg6sXnZIgYrOxWGvbx+QMq
mNRpvQDCLVzJN0SgVdjfqAG2TG71dX2AjcX9EQujGOHFudUY4xl0Sl082yY8iA5a
+HS3atS/ZKqvuLS1gkmiWam8Kr4QLm6BIQ+4s2mC9Vbt3WDE5UDEpNyF9RNU6e4l
WCyhpFggNRMadZNcf8ifbN3b+f60jM0NnpgJ3Bm6BGyECXO8blhGMea/qP1xrL8o
Fwrdw5lEPSror5UquAsVF/D1B8m0zYroLkakHJroXpdlVskGr2SvB9AWu0qjI4S4
yYeth4Mwn6uzNSOFzeH+anlvDfmliH6NmCYQvAi4/t/ObgDMtnjwcasgAH/s2yF1
3c13dstyqeL73nH9tRUx1QwqNPVDnD8vLxyLRoPcD0yMhlyoG/spf009GALQJa6p
MOhnqLl+jZTwIRqHMD3+oaZbovLFUl8borlA3VuQODsLmzoRr9ftwiUgHOieStaK
15R9jnP73lVDYmF6X1rBZQnxh2Xv7fNs6iIsow+7msvqYjgvZ91/OH69PR7Dw8/b
H02fsQtziytVd/wLOccrxkn/JExnIoSN3Eji+HnfhfFnnCndW8Pkf5EkY1sVLJe/
68aVWLRtQ0wsbIA2C/F5IWa/x9BHp9K0sxlPTq6cBouUZyWFZTIW2CW4YYa3qRIp
F9MvyIWp2+lynJ+3BfBxfkFVpPpvVKu5/RGsPBCNUgcxgBu8SYzIBnbcVyzXhcNn
9nCVsrf94Sj86uVoVglsXx5O1hAY28G0MZkiWpOK+1304Ks3gCi8KmQ33PjYJjj9
kpC/pegVN2yLVF2ablpJaLvtXBIc5Oxy/WlOs/t1jtgpyGvXYpx8DYd28uC0zwTg
n0eZhGfQvyq1EtJjZRmBgFgnDRMQQIw+gCVpcY1QHrPHqxVib1XnnuHeu39KwRoU
RpiEhkkOeK/B89Z6xi8mGwsG6Zbfyf7bJbKaRZEFrcOvmgsFvO5fz9V0ULgpje4M
eM+zGBzzCcf/Qn76rnXxd/lVk2r8DRMQNfTvUuWT82iM+zwlEyoKk3AEyPpJT5dU
OBnPy8THuLpnq2W0HylC9OBuMY7SOQJfyztVy7CraTsFnH5RXPqUdZpZ4mZ8w5+m
0i6NvCL+hEh8EjyYRf7LAIvabNsAnTuykINhH10RUhK06G3D4DWtXF/up6149W3T
yUBTETBLCXfSV7svOPfoTdek8tEtL4cFpQ1JszqWsCxoJkGMY/SI/n2Scl4zMNoZ
leEzxqlWEf4Ugrm9uFi0U8Tgc4HobneFTfO6RnlxnhxV5rIKknaXvnHW9M9BneW3
iRk7Hksd5L1HfqqBJ/ybQTD47BHZ0Bi6km+d232dNabscAhOzVvdQskY0tJqVyKO
Kf7CXhCyMwKNnNx+1nH+WQ==
//pragma protect end_data_block
//pragma protect digest_block
W/z2334kvpnA6+eEw1UKoV9h/tw=
//pragma protect end_digest_block
//pragma protect end_protected
