module CHIP(
            clk,
            rst_n,
            IN_VALID,
            MODE,
            FFT2D_IN_R,
            FFT2D_IN_I,
            OUT_VALID,
            FFT2D_OUT_R,
            FFT2D_OUT_I
);
input         clk, rst_n, IN_VALID, MODE;
input  [18:0] FFT2D_IN_R, FFT2D_IN_I;

output        OUT_VALID;
output [18:0] FFT2D_OUT_R, FFT2D_OUT_I;


wire        C_clk, C_rst_n, C_IN_VALID, C_MODE;
wire [18:0] C_FFT2D_IN_R, C_FFT2D_IN_I;

wire        C_OUT_VALID;
wire [18:0] C_FFT2D_OUT_R, C_FFT2D_OUT_I;

wire BUF_clk;
CLKBUFX20 buf0(.A(C_clk),.Y(BUF_clk));

FFT2D u_FFT2D(
    .clk(BUF_clk),
    .rst_n(C_rst_n),
    .IN_VALID(C_IN_VALID),
    .MODE(C_MODE),
    .FFT2D_IN_R(C_FFT2D_IN_R),
    .FFT2D_IN_I(C_FFT2D_IN_I),
    .OUT_VALID(C_OUT_VALID),
    .FFT2D_OUT_R(C_FFT2D_OUT_R),
    .FFT2D_OUT_I(C_FFT2D_OUT_I)
    );

// Input Pads
P8C I_CLK      ( .Y(C_clk),        .P(clk),        .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b0), .CSEN(1'b1) );
P8C I_RESET    ( .Y(C_rst_n),      .P(rst_n),      .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_VALID    ( .Y(C_IN_VALID),   .P(IN_VALID),   .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );

P4C I_MODE     ( .Y(C_MODE), .P(MODE), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );

P4C I_FFT2D_IN_R_0     ( .Y(C_FFT2D_IN_R[0]), .P(FFT2D_IN_R[0]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_FFT2D_IN_R_1     ( .Y(C_FFT2D_IN_R[1]), .P(FFT2D_IN_R[1]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_FFT2D_IN_R_2     ( .Y(C_FFT2D_IN_R[2]), .P(FFT2D_IN_R[2]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_FFT2D_IN_R_3     ( .Y(C_FFT2D_IN_R[3]), .P(FFT2D_IN_R[3]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_FFT2D_IN_R_4     ( .Y(C_FFT2D_IN_R[4]), .P(FFT2D_IN_R[4]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_FFT2D_IN_R_5     ( .Y(C_FFT2D_IN_R[5]), .P(FFT2D_IN_R[5]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_FFT2D_IN_R_6     ( .Y(C_FFT2D_IN_R[6]), .P(FFT2D_IN_R[6]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_FFT2D_IN_R_7     ( .Y(C_FFT2D_IN_R[7]), .P(FFT2D_IN_R[7]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_FFT2D_IN_R_8     ( .Y(C_FFT2D_IN_R[8]), .P(FFT2D_IN_R[8]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_FFT2D_IN_R_9     ( .Y(C_FFT2D_IN_R[9]), .P(FFT2D_IN_R[9]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_FFT2D_IN_R_10     ( .Y(C_FFT2D_IN_R[10]), .P(FFT2D_IN_R[10]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_FFT2D_IN_R_11     ( .Y(C_FFT2D_IN_R[11]), .P(FFT2D_IN_R[11]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_FFT2D_IN_R_12     ( .Y(C_FFT2D_IN_R[12]), .P(FFT2D_IN_R[12]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_FFT2D_IN_R_13     ( .Y(C_FFT2D_IN_R[13]), .P(FFT2D_IN_R[13]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_FFT2D_IN_R_14     ( .Y(C_FFT2D_IN_R[14]), .P(FFT2D_IN_R[14]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_FFT2D_IN_R_15     ( .Y(C_FFT2D_IN_R[15]), .P(FFT2D_IN_R[15]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_FFT2D_IN_R_16     ( .Y(C_FFT2D_IN_R[16]), .P(FFT2D_IN_R[16]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_FFT2D_IN_R_17     ( .Y(C_FFT2D_IN_R[17]), .P(FFT2D_IN_R[17]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_FFT2D_IN_R_18     ( .Y(C_FFT2D_IN_R[18]), .P(FFT2D_IN_R[18]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );

P4C I_FFT2D_IN_I_0     ( .Y(C_FFT2D_IN_I[0]), .P(FFT2D_IN_I[0]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_FFT2D_IN_I_1     ( .Y(C_FFT2D_IN_I[1]), .P(FFT2D_IN_I[1]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_FFT2D_IN_I_2     ( .Y(C_FFT2D_IN_I[2]), .P(FFT2D_IN_I[2]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_FFT2D_IN_I_3     ( .Y(C_FFT2D_IN_I[3]), .P(FFT2D_IN_I[3]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_FFT2D_IN_I_4     ( .Y(C_FFT2D_IN_I[4]), .P(FFT2D_IN_I[4]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_FFT2D_IN_I_5     ( .Y(C_FFT2D_IN_I[5]), .P(FFT2D_IN_I[5]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_FFT2D_IN_I_6     ( .Y(C_FFT2D_IN_I[6]), .P(FFT2D_IN_I[6]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_FFT2D_IN_I_7     ( .Y(C_FFT2D_IN_I[7]), .P(FFT2D_IN_I[7]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_FFT2D_IN_I_8     ( .Y(C_FFT2D_IN_I[8]), .P(FFT2D_IN_I[8]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_FFT2D_IN_I_9     ( .Y(C_FFT2D_IN_I[9]), .P(FFT2D_IN_I[9]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_FFT2D_IN_I_10     ( .Y(C_FFT2D_IN_I[10]), .P(FFT2D_IN_I[10]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_FFT2D_IN_I_11     ( .Y(C_FFT2D_IN_I[11]), .P(FFT2D_IN_I[11]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_FFT2D_IN_I_12     ( .Y(C_FFT2D_IN_I[12]), .P(FFT2D_IN_I[12]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_FFT2D_IN_I_13     ( .Y(C_FFT2D_IN_I[13]), .P(FFT2D_IN_I[13]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_FFT2D_IN_I_14     ( .Y(C_FFT2D_IN_I[14]), .P(FFT2D_IN_I[14]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_FFT2D_IN_I_15     ( .Y(C_FFT2D_IN_I[15]), .P(FFT2D_IN_I[15]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_FFT2D_IN_I_16     ( .Y(C_FFT2D_IN_I[16]), .P(FFT2D_IN_I[16]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_FFT2D_IN_I_17     ( .Y(C_FFT2D_IN_I[17]), .P(FFT2D_IN_I[17]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_FFT2D_IN_I_18     ( .Y(C_FFT2D_IN_I[18]), .P(FFT2D_IN_I[18]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );

// Output Pads
P8C O_VALID    ( .A(C_OUT_VALID),   .P(OUT_VALID), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );

P8C O_FFT2D_OUT_R_0     ( .A(C_FFT2D_OUT_R[0]), .P(FFT2D_OUT_R[0]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P8C O_FFT2D_OUT_R_1     ( .A(C_FFT2D_OUT_R[1]), .P(FFT2D_OUT_R[1]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P8C O_FFT2D_OUT_R_2     ( .A(C_FFT2D_OUT_R[2]), .P(FFT2D_OUT_R[2]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P8C O_FFT2D_OUT_R_3     ( .A(C_FFT2D_OUT_R[3]), .P(FFT2D_OUT_R[3]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P8C O_FFT2D_OUT_R_4     ( .A(C_FFT2D_OUT_R[4]), .P(FFT2D_OUT_R[4]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P8C O_FFT2D_OUT_R_5     ( .A(C_FFT2D_OUT_R[5]), .P(FFT2D_OUT_R[5]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P8C O_FFT2D_OUT_R_6     ( .A(C_FFT2D_OUT_R[6]), .P(FFT2D_OUT_R[6]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P8C O_FFT2D_OUT_R_7     ( .A(C_FFT2D_OUT_R[7]), .P(FFT2D_OUT_R[7]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P8C O_FFT2D_OUT_R_8     ( .A(C_FFT2D_OUT_R[8]), .P(FFT2D_OUT_R[8]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P8C O_FFT2D_OUT_R_9     ( .A(C_FFT2D_OUT_R[9]), .P(FFT2D_OUT_R[9]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P8C O_FFT2D_OUT_R_10     ( .A(C_FFT2D_OUT_R[10]), .P(FFT2D_OUT_R[10]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P8C O_FFT2D_OUT_R_11     ( .A(C_FFT2D_OUT_R[11]), .P(FFT2D_OUT_R[11]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P8C O_FFT2D_OUT_R_12     ( .A(C_FFT2D_OUT_R[12]), .P(FFT2D_OUT_R[12]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P8C O_FFT2D_OUT_R_13     ( .A(C_FFT2D_OUT_R[13]), .P(FFT2D_OUT_R[13]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P8C O_FFT2D_OUT_R_14     ( .A(C_FFT2D_OUT_R[14]), .P(FFT2D_OUT_R[14]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P8C O_FFT2D_OUT_R_15     ( .A(C_FFT2D_OUT_R[15]), .P(FFT2D_OUT_R[15]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P8C O_FFT2D_OUT_R_16     ( .A(C_FFT2D_OUT_R[16]), .P(FFT2D_OUT_R[16]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P8C O_FFT2D_OUT_R_17     ( .A(C_FFT2D_OUT_R[17]), .P(FFT2D_OUT_R[17]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P8C O_FFT2D_OUT_R_18     ( .A(C_FFT2D_OUT_R[18]), .P(FFT2D_OUT_R[18]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );

P8C O_FFT2D_OUT_I_0     ( .A(C_FFT2D_OUT_I[0]), .P(FFT2D_OUT_I[0]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P8C O_FFT2D_OUT_I_1     ( .A(C_FFT2D_OUT_I[1]), .P(FFT2D_OUT_I[1]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P8C O_FFT2D_OUT_I_2     ( .A(C_FFT2D_OUT_I[2]), .P(FFT2D_OUT_I[2]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P8C O_FFT2D_OUT_I_3     ( .A(C_FFT2D_OUT_I[3]), .P(FFT2D_OUT_I[3]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P8C O_FFT2D_OUT_I_4     ( .A(C_FFT2D_OUT_I[4]), .P(FFT2D_OUT_I[4]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P8C O_FFT2D_OUT_I_5     ( .A(C_FFT2D_OUT_I[5]), .P(FFT2D_OUT_I[5]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P8C O_FFT2D_OUT_I_6     ( .A(C_FFT2D_OUT_I[6]), .P(FFT2D_OUT_I[6]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P8C O_FFT2D_OUT_I_7     ( .A(C_FFT2D_OUT_I[7]), .P(FFT2D_OUT_I[7]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P8C O_FFT2D_OUT_I_8     ( .A(C_FFT2D_OUT_I[8]), .P(FFT2D_OUT_I[8]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P8C O_FFT2D_OUT_I_9     ( .A(C_FFT2D_OUT_I[9]), .P(FFT2D_OUT_I[9]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P8C O_FFT2D_OUT_I_10     ( .A(C_FFT2D_OUT_I[10]), .P(FFT2D_OUT_I[10]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P8C O_FFT2D_OUT_I_11     ( .A(C_FFT2D_OUT_I[11]), .P(FFT2D_OUT_I[11]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P8C O_FFT2D_OUT_I_12     ( .A(C_FFT2D_OUT_I[12]), .P(FFT2D_OUT_I[12]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P8C O_FFT2D_OUT_I_13     ( .A(C_FFT2D_OUT_I[13]), .P(FFT2D_OUT_I[13]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P8C O_FFT2D_OUT_I_14     ( .A(C_FFT2D_OUT_I[14]), .P(FFT2D_OUT_I[14]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P8C O_FFT2D_OUT_I_15     ( .A(C_FFT2D_OUT_I[15]), .P(FFT2D_OUT_I[15]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P8C O_FFT2D_OUT_I_16     ( .A(C_FFT2D_OUT_I[16]), .P(FFT2D_OUT_I[16]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P8C O_FFT2D_OUT_I_17     ( .A(C_FFT2D_OUT_I[17]), .P(FFT2D_OUT_I[17]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P8C O_FFT2D_OUT_I_18     ( .A(C_FFT2D_OUT_I[18]), .P(FFT2D_OUT_I[18]), .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );

//I/O power 3.3V pads  (DVDD + DGND) at least 8 pairs
PVDDR VDDP0 ();
PVSSR GNDP0 ();
PVDDR VDDP1 ();
PVSSR GNDP1 ();
PVDDR VDDP2 ();
PVSSR GNDP2 ();
PVDDR VDDP3 ();
PVSSR GNDP3 ();
PVDDR VDDP4 ();
PVSSR GNDP4 ();
PVDDR VDDP5 ();
PVSSR GNDP5 ();
PVDDR VDDP6 ();
PVSSR GNDP6 ();
PVDDR VDDP7 ();
PVSSR GNDP7 ();

//Core poweri 1.8V pads  (VDD + GND) at least 2 pairs, (don't placed near the corner).
PVDDC VDDC0 ();
PVSSC GNDC0 ();
PVDDC VDDC1 ();
PVSSC GNDC1 ();

endmodule
/////////////////////////////////////////////////////////////
// Created by: Synopsys DC Ultra(TM) in wire load mode
// Version   : K-2015.06-SP1
// Date      : Wed Jan 16 19:10:13 2019
/////////////////////////////////////////////////////////////


module FFT2D ( clk, rst_n, IN_VALID, MODE, FFT2D_IN_R, FFT2D_IN_I, OUT_VALID, 
        FFT2D_OUT_R, FFT2D_OUT_I );
  input [18:0] FFT2D_IN_R;
  input [18:0] FFT2D_IN_I;
  output [18:0] FFT2D_OUT_R;
  output [18:0] FFT2D_OUT_I;
  input clk, rst_n, IN_VALID, MODE;
  output OUT_VALID;
  wire   WEN, is_row, mode_val, N1156, N1157, N1158, N1159, N1160, N1161,
         N1162, N1163, N1164, N1165, N1166, N1236, N1237, N1238, N1239, N1240,
         N1241, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567,
         DP_OP_132J1_122_4436_n2999, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2846, n2847,
         n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
         n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
         n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3268, n3269,
         n3270, n3271, n3272, n3273, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
         n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
         n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678;
  wire   [10:0] A;
  wire   [3:0] cs;
  wire   [5:0] lay_cnt;
  wire   [4:0] sequence_cnt;
  wire   [10:0] in_out_cnt;
  wire   [18:0] D_real;
  wire   [18:0] D_imag;
  wire   [17:0] butt_a_real;
  wire   [18:0] butt_a_imag;
  wire   [18:0] butt_b_real;
  wire   [18:0] butt_b_imag;
  tri   [37:0] Q;

  RA1SH1 SRAM_mem ( .Q(Q), .A(A), .D({D_real, D_imag}), .CLK(clk), .CEN(1'b0), 
        .OEN(1'b0), .WEN(WEN) );
  DFFRHQX4 cs_reg_0_ ( .D(n564), .CK(clk), .RN(rst_n), .Q(cs[0]) );
  DFFRHQXL is_row_reg ( .D(n558), .CK(clk), .RN(rst_n), .Q(is_row) );
  DFFRHQX4 cs_reg_1_ ( .D(n565), .CK(clk), .RN(rst_n), .Q(cs[1]) );
  DFFRHQX4 cs_reg_2_ ( .D(n566), .CK(clk), .RN(rst_n), .Q(cs[2]) );
  DFFRHQXL in_out_cnt_reg_0_ ( .D(N1156), .CK(clk), .RN(rst_n), .Q(
        in_out_cnt[0]) );
  DFFRHQXL in_out_cnt_reg_1_ ( .D(N1157), .CK(clk), .RN(rst_n), .Q(
        in_out_cnt[1]) );
  DFFRHQXL in_out_cnt_reg_2_ ( .D(N1158), .CK(clk), .RN(rst_n), .Q(
        in_out_cnt[2]) );
  DFFRHQXL in_out_cnt_reg_3_ ( .D(N1159), .CK(clk), .RN(rst_n), .Q(
        in_out_cnt[3]) );
  DFFRHQXL in_out_cnt_reg_4_ ( .D(N1160), .CK(clk), .RN(rst_n), .Q(
        in_out_cnt[4]) );
  DFFRHQXL in_out_cnt_reg_5_ ( .D(N1161), .CK(clk), .RN(rst_n), .Q(
        in_out_cnt[5]) );
  DFFRHQXL in_out_cnt_reg_6_ ( .D(N1162), .CK(clk), .RN(rst_n), .Q(
        in_out_cnt[6]) );
  DFFRHQXL in_out_cnt_reg_7_ ( .D(N1163), .CK(clk), .RN(rst_n), .Q(
        in_out_cnt[7]) );
  DFFRHQXL in_out_cnt_reg_8_ ( .D(N1164), .CK(clk), .RN(rst_n), .Q(
        in_out_cnt[8]) );
  DFFRHQXL in_out_cnt_reg_9_ ( .D(N1165), .CK(clk), .RN(rst_n), .Q(
        in_out_cnt[9]) );
  DFFRHQXL in_out_cnt_reg_10_ ( .D(N1166), .CK(clk), .RN(rst_n), .Q(
        in_out_cnt[10]) );
  DFFRHQX4 cs_reg_3_ ( .D(n567), .CK(clk), .RN(rst_n), .Q(cs[3]) );
  DFFRHQXL lay_cnt_reg_1_ ( .D(N1237), .CK(clk), .RN(rst_n), .Q(lay_cnt[1]) );
  DFFRHQX4 lay_cnt_reg_2_ ( .D(N1238), .CK(clk), .RN(rst_n), .Q(lay_cnt[2]) );
  DFFRHQX4 lay_cnt_reg_3_ ( .D(N1239), .CK(clk), .RN(rst_n), .Q(lay_cnt[3]) );
  DFFRHQX2 lay_cnt_reg_5_ ( .D(N1241), .CK(clk), .RN(rst_n), .Q(lay_cnt[5]) );
  DFFRHQXL mode_val_reg ( .D(n557), .CK(clk), .RN(rst_n), .Q(mode_val) );
  DFFRHQX4 butt_b_imag_reg_9_ ( .D(n556), .CK(clk), .RN(rst_n), .Q(
        butt_b_imag[9]) );
  DFFRHQX4 butt_b_imag_reg_6_ ( .D(n550), .CK(clk), .RN(rst_n), .Q(
        butt_b_imag[6]) );
  DFFRHQX4 butt_b_imag_reg_4_ ( .D(n546), .CK(clk), .RN(rst_n), .Q(
        butt_b_imag[4]) );
  DFFRHQX4 butt_a_imag_reg_4_ ( .D(n545), .CK(clk), .RN(rst_n), .Q(
        butt_a_imag[4]) );
  DFFRHQX4 butt_b_real_reg_16_ ( .D(n538), .CK(clk), .RN(rst_n), .Q(
        butt_b_real[16]) );
  DFFRHQX4 butt_a_real_reg_16_ ( .D(n537), .CK(clk), .RN(rst_n), .Q(
        butt_a_real[16]) );
  DFFRHQX4 butt_a_real_reg_14_ ( .D(n533), .CK(clk), .RN(rst_n), .Q(
        butt_a_real[14]) );
  DFFRHQX4 butt_a_real_reg_11_ ( .D(n527), .CK(clk), .RN(rst_n), .Q(
        butt_a_real[11]) );
  DFFRHQX4 butt_b_imag_reg_2_ ( .D(n526), .CK(clk), .RN(rst_n), .Q(
        butt_b_imag[2]) );
  DFFRHQX4 butt_b_real_reg_10_ ( .D(n524), .CK(clk), .RN(rst_n), .Q(
        butt_b_real[10]) );
  DFFRHQX4 butt_a_real_reg_10_ ( .D(n523), .CK(clk), .RN(rst_n), .Q(
        butt_a_real[10]) );
  DFFRHQX4 butt_b_real_reg_8_ ( .D(n520), .CK(clk), .RN(rst_n), .Q(
        butt_b_real[8]) );
  DFFRHQX4 butt_a_real_reg_8_ ( .D(n519), .CK(clk), .RN(rst_n), .Q(
        butt_a_real[8]) );
  DFFRHQX4 butt_a_real_reg_6_ ( .D(n515), .CK(clk), .RN(rst_n), .Q(
        butt_a_real[6]) );
  DFFRHQX4 butt_b_real_reg_5_ ( .D(n514), .CK(clk), .RN(rst_n), .Q(
        butt_b_real[5]) );
  DFFRHQX4 butt_a_real_reg_5_ ( .D(n513), .CK(clk), .RN(rst_n), .Q(
        butt_a_real[5]) );
  DFFRHQX4 butt_a_real_reg_4_ ( .D(n511), .CK(clk), .RN(rst_n), .Q(
        butt_a_real[4]) );
  DFFRHQX4 butt_a_real_reg_2_ ( .D(n507), .CK(clk), .RN(rst_n), .Q(
        butt_a_real[2]) );
  DFFRHQX2 butt_b_real_reg_1_ ( .D(n506), .CK(clk), .RN(rst_n), .Q(
        butt_b_real[1]) );
  DFFRHQX4 butt_a_imag_reg_16_ ( .D(n495), .CK(clk), .RN(rst_n), .Q(
        butt_a_imag[16]) );
  DFFRHQX4 butt_b_imag_reg_12_ ( .D(n488), .CK(clk), .RN(rst_n), .Q(
        butt_b_imag[12]) );
  DFFRHQX4 butt_a_imag_reg_12_ ( .D(n487), .CK(clk), .RN(rst_n), .Q(
        butt_a_imag[12]) );
  DFFRHQX4 butt_a_imag_reg_11_ ( .D(n485), .CK(clk), .RN(rst_n), .Q(
        butt_a_imag[11]) );
  DFFRHQX4 butt_b_imag_reg_10_ ( .D(n484), .CK(clk), .RN(rst_n), .Q(
        butt_b_imag[10]) );
  DFFRHQX2 butt_a_imag_reg_0_ ( .D(n481), .CK(clk), .RN(rst_n), .Q(
        butt_a_imag[0]) );
  DFFRHQX4 butt_a_imag_reg_10_ ( .D(n483), .CK(clk), .RN(rst_n), .Q(
        butt_a_imag[10]) );
  DFFRHQX4 butt_b_real_reg_6_ ( .D(n516), .CK(clk), .RN(rst_n), .Q(
        butt_b_real[6]) );
  DFFRHQX4 butt_a_imag_reg_5_ ( .D(n547), .CK(clk), .RN(rst_n), .Q(
        butt_a_imag[5]) );
  DFFRHQX4 butt_a_real_reg_3_ ( .D(n509), .CK(clk), .RN(rst_n), .Q(
        butt_a_real[3]) );
  DFFRHQX4 butt_a_real_reg_7_ ( .D(n517), .CK(clk), .RN(rst_n), .Q(
        butt_a_real[7]) );
  DFFRHQX4 butt_a_imag_reg_13_ ( .D(n489), .CK(clk), .RN(rst_n), .Q(
        butt_a_imag[13]) );
  DFFRHQX4 butt_a_imag_reg_3_ ( .D(n543), .CK(clk), .RN(rst_n), .Q(
        butt_a_imag[3]) );
  DFFRHQX4 butt_b_real_reg_3_ ( .D(n510), .CK(clk), .RN(rst_n), .Q(
        butt_b_real[3]) );
  DFFRHQX4 lay_cnt_reg_4_ ( .D(N1240), .CK(clk), .RN(rst_n), .Q(lay_cnt[4]) );
  DFFRHQX4 butt_b_real_reg_2_ ( .D(n508), .CK(clk), .RN(rst_n), .Q(
        butt_b_real[2]) );
  DFFRHQX4 butt_a_real_reg_9_ ( .D(n521), .CK(clk), .RN(rst_n), .Q(
        butt_a_real[9]) );
  DFFRHQX4 butt_b_real_reg_7_ ( .D(n518), .CK(clk), .RN(rst_n), .Q(
        butt_b_real[7]) );
  DFFSX1 OUT_VALID_reg ( .D(n4675), .CK(clk), .SN(rst_n), .QN(OUT_VALID) );
  DFFSX1 sequence_cnt_reg_1_ ( .D(n562), .CK(clk), .SN(rst_n), .Q(
        sequence_cnt[1]), .QN(n4678) );
  DFFSX1 sequence_cnt_reg_0_ ( .D(n563), .CK(clk), .SN(rst_n), .Q(
        sequence_cnt[0]) );
  DFFSX1 sequence_cnt_reg_4_ ( .D(n559), .CK(clk), .SN(rst_n), .Q(
        sequence_cnt[4]) );
  DFFSX1 sequence_cnt_reg_3_ ( .D(n560), .CK(clk), .SN(rst_n), .Q(
        sequence_cnt[3]) );
  DFFSX1 sequence_cnt_reg_2_ ( .D(n561), .CK(clk), .SN(rst_n), .Q(
        sequence_cnt[2]), .QN(n4676) );
  DFFRX1 lay_cnt_reg_0_ ( .D(N1236), .CK(clk), .RN(rst_n), .Q(lay_cnt[0]), 
        .QN(n4677) );
  DFFSHQX4 butt_a_imag_reg_1_ ( .D(n4670), .CK(clk), .SN(rst_n), .Q(n4671) );
  DFFRHQX4 butt_a_imag_reg_15_ ( .D(n493), .CK(clk), .RN(rst_n), .Q(
        butt_a_imag[15]) );
  DFFRHQX4 butt_b_imag_reg_13_ ( .D(n490), .CK(clk), .RN(rst_n), .Q(
        butt_b_imag[13]) );
  DFFRHQX4 butt_a_real_reg_15_ ( .D(n535), .CK(clk), .RN(rst_n), .Q(
        butt_a_real[15]) );
  DFFRHQX1 butt_b_imag_reg_0_ ( .D(n482), .CK(clk), .RN(rst_n), .Q(
        butt_b_imag[0]) );
  DFFRHQX2 butt_b_real_reg_13_ ( .D(n532), .CK(clk), .RN(rst_n), .Q(
        butt_b_real[13]) );
  DFFRHQX2 butt_a_imag_reg_18_ ( .D(n499), .CK(clk), .RN(rst_n), .Q(
        butt_a_imag[18]) );
  DFFRHQX2 butt_a_imag_reg_7_ ( .D(n551), .CK(clk), .RN(rst_n), .Q(
        butt_a_imag[7]) );
  DFFRHQX2 butt_a_imag_reg_8_ ( .D(n553), .CK(clk), .RN(rst_n), .Q(
        butt_a_imag[8]) );
  DFFRHQX2 butt_b_imag_reg_14_ ( .D(n492), .CK(clk), .RN(rst_n), .Q(
        butt_b_imag[14]) );
  DFFRHQX2 butt_b_real_reg_14_ ( .D(n534), .CK(clk), .RN(rst_n), .Q(
        butt_b_real[14]) );
  DFFRHQX2 butt_b_imag_reg_16_ ( .D(n496), .CK(clk), .RN(rst_n), .Q(
        butt_b_imag[16]) );
  DFFRHQX2 butt_b_imag_reg_1_ ( .D(n504), .CK(clk), .RN(rst_n), .Q(
        butt_b_imag[1]) );
  DFFRHQX2 butt_a_real_reg_13_ ( .D(n531), .CK(clk), .RN(rst_n), .Q(
        butt_a_real[13]) );
  DFFRHQX2 butt_b_imag_reg_15_ ( .D(n494), .CK(clk), .RN(rst_n), .Q(
        butt_b_imag[15]) );
  DFFRHQX2 butt_a_imag_reg_14_ ( .D(n491), .CK(clk), .RN(rst_n), .Q(
        butt_a_imag[14]) );
  DFFRHQX2 butt_b_real_reg_15_ ( .D(n536), .CK(clk), .RN(rst_n), .Q(
        butt_b_real[15]) );
  DFFRHQX1 butt_b_imag_reg_8_ ( .D(n554), .CK(clk), .RN(rst_n), .Q(
        butt_b_imag[8]) );
  DFFRHQX2 butt_b_real_reg_17_ ( .D(n540), .CK(clk), .RN(rst_n), .Q(
        butt_b_real[17]) );
  DFFRHQX2 butt_b_real_reg_12_ ( .D(n530), .CK(clk), .RN(rst_n), .Q(
        butt_b_real[12]) );
  DFFRHQX2 butt_b_real_reg_11_ ( .D(n528), .CK(clk), .RN(rst_n), .Q(
        butt_b_real[11]) );
  DFFRHQX2 butt_b_real_reg_4_ ( .D(n512), .CK(clk), .RN(rst_n), .Q(
        butt_b_real[4]) );
  DFFRHQX2 butt_a_real_reg_12_ ( .D(n529), .CK(clk), .RN(rst_n), .Q(
        butt_a_real[12]) );
  DFFRHQX2 butt_a_imag_reg_6_ ( .D(n549), .CK(clk), .RN(rst_n), .Q(
        butt_a_imag[6]) );
  DFFRHQX1 butt_b_imag_reg_3_ ( .D(n544), .CK(clk), .RN(rst_n), .Q(
        butt_b_imag[3]) );
  DFFRHQX2 butt_b_real_reg_9_ ( .D(n522), .CK(clk), .RN(rst_n), .Q(
        butt_b_real[9]) );
  DFFRHQX2 butt_b_real_reg_18_ ( .D(n542), .CK(clk), .RN(rst_n), .Q(
        butt_b_real[18]) );
  DFFRHQX2 butt_b_imag_reg_17_ ( .D(n498), .CK(clk), .RN(rst_n), .Q(
        butt_b_imag[17]) );
  DFFRHQX2 butt_a_imag_reg_17_ ( .D(n497), .CK(clk), .RN(rst_n), .Q(
        butt_a_imag[17]) );
  DFFRHQX2 butt_b_imag_reg_7_ ( .D(n552), .CK(clk), .RN(rst_n), .Q(
        butt_b_imag[7]) );
  DFFRHQX2 butt_a_real_reg_17_ ( .D(n539), .CK(clk), .RN(rst_n), .Q(
        butt_a_real[17]) );
  DFFSHQX2 butt_a_real_reg_18_ ( .D(n4672), .CK(clk), .SN(rst_n), .Q(n4673) );
  DFFRHQX2 butt_a_imag_reg_2_ ( .D(n525), .CK(clk), .RN(rst_n), .Q(
        butt_a_imag[2]) );
  DFFRHQX2 butt_a_imag_reg_9_ ( .D(n555), .CK(clk), .RN(rst_n), .Q(
        butt_a_imag[9]) );
  DFFRHQX2 butt_a_real_reg_1_ ( .D(n505), .CK(clk), .RN(rst_n), .Q(
        butt_a_real[1]) );
  DFFRHQX2 butt_b_imag_reg_11_ ( .D(n486), .CK(clk), .RN(rst_n), .Q(
        butt_b_imag[11]) );
  DFFRHQX2 butt_b_imag_reg_5_ ( .D(n548), .CK(clk), .RN(rst_n), .Q(
        butt_b_imag[5]) );
  DFFSX1 butt_b_real_reg_0_ ( .D(n4674), .CK(clk), .SN(rst_n), .Q(
        DP_OP_132J1_122_4436_n2999), .QN(butt_b_real[0]) );
  DFFRHQX2 butt_b_imag_reg_18_ ( .D(n500), .CK(clk), .RN(rst_n), .Q(
        butt_b_imag[18]) );
  DFFRHQX1 butt_a_real_reg_0_ ( .D(n501), .CK(clk), .RN(rst_n), .Q(
        butt_a_real[0]) );
  NOR2X1 U696 ( .A(in_out_cnt[0]), .B(n4664), .Y(N1156) );
  NOR2X1 U697 ( .A(n4102), .B(n3763), .Y(N1238) );
  NOR2X1 U698 ( .A(sequence_cnt[4]), .B(n3758), .Y(n3761) );
  NOR2X1 U699 ( .A(n1123), .B(n4592), .Y(n4306) );
  INVX2 U700 ( .A(n619), .Y(n620) );
  NOR2X1 U701 ( .A(n4352), .B(n4563), .Y(n4358) );
  NAND2X1 U702 ( .A(n4111), .B(n4675), .Y(n4661) );
  XOR2X2 U703 ( .A(n2331), .B(n1115), .Y(n1090) );
  NAND2X1 U704 ( .A(n834), .B(n3573), .Y(n833) );
  NAND3X2 U705 ( .A(rst_n), .B(OUT_VALID), .C(n3858), .Y(n3866) );
  NOR2X1 U706 ( .A(n3858), .B(n3857), .Y(n3859) );
  NAND2X2 U707 ( .A(n803), .B(n3548), .Y(n802) );
  XOR2X2 U708 ( .A(n854), .B(n659), .Y(n4433) );
  NOR2X1 U709 ( .A(lay_cnt[1]), .B(is_row), .Y(n4623) );
  AND2X1 U710 ( .A(n4028), .B(n3999), .Y(n658) );
  NOR2X1 U711 ( .A(n3821), .B(lay_cnt[1]), .Y(n4650) );
  CLKINVX2 U712 ( .A(n914), .Y(n803) );
  NOR2X1 U713 ( .A(n4030), .B(n4033), .Y(n4037) );
  NOR2X1 U714 ( .A(n3567), .B(n3570), .Y(n3568) );
  NAND2X1 U715 ( .A(n4111), .B(n3762), .Y(n2371) );
  NOR2X1 U716 ( .A(n3772), .B(n3840), .Y(n3771) );
  NOR2X1 U717 ( .A(n4644), .B(mode_val), .Y(n2056) );
  NOR2X1 U718 ( .A(n3833), .B(n4657), .Y(n4663) );
  NOR2X1 U719 ( .A(n605), .B(n3811), .Y(n3780) );
  NAND2X2 U720 ( .A(n2372), .B(n2277), .Y(n4024) );
  OR2X1 U721 ( .A(n3523), .B(n3522), .Y(n3521) );
  NOR2X2 U722 ( .A(n3692), .B(n3688), .Y(n2372) );
  NAND2X1 U723 ( .A(n2282), .B(n2281), .Y(n4004) );
  NOR2X2 U724 ( .A(n3425), .B(n3426), .Y(n4463) );
  NAND2X2 U725 ( .A(n2337), .B(n2342), .Y(n2345) );
  NOR2X2 U726 ( .A(n4104), .B(lay_cnt[0]), .Y(n4184) );
  INVX2 U727 ( .A(IN_VALID), .Y(n4111) );
  NAND2X1 U728 ( .A(n3395), .B(n3394), .Y(n3408) );
  NAND2X2 U729 ( .A(n902), .B(n703), .Y(n4472) );
  NOR2X1 U730 ( .A(n962), .B(n963), .Y(n2343) );
  NOR2X1 U731 ( .A(n1461), .B(n1460), .Y(n4416) );
  NOR2X1 U732 ( .A(n1624), .B(n1623), .Y(n3932) );
  OR2XL U733 ( .A(n1850), .B(n1851), .Y(n1854) );
  OR2XL U734 ( .A(n2153), .B(n2154), .Y(n2157) );
  NOR2X1 U735 ( .A(n3322), .B(n3321), .Y(n4292) );
  INVX2 U736 ( .A(n1931), .Y(n788) );
  OR2XL U737 ( .A(n1448), .B(n1447), .Y(n1450) );
  OAI2BB1X2 U738 ( .A0N(n1021), .A1N(n3371), .B0(n3354), .Y(n3379) );
  OAI2BB1X2 U739 ( .A0N(n1732), .A1N(n694), .B0(n693), .Y(n1853) );
  NAND2X1 U740 ( .A(n905), .B(n904), .Y(n1855) );
  ADDFX1 U741 ( .A(n1457), .B(n1456), .CI(n1455), .CO(n1458), .S(n1448) );
  OR2XL U742 ( .A(n2600), .B(n2599), .Y(n2525) );
  INVX2 U743 ( .A(n1818), .Y(n1856) );
  ADDFX2 U744 ( .A(n1437), .B(n1436), .CI(n1435), .CO(n1457), .S(n1430) );
  ADDFHX1 U745 ( .A(n2876), .B(n2875), .CI(n2874), .CO(n2946), .S(n3356) );
  ADDFHX1 U746 ( .A(n1587), .B(n1585), .CI(n1586), .CO(n1696), .S(n1617) );
  XNOR3X2 U747 ( .A(n2810), .B(n1050), .C(n2809), .Y(n2951) );
  NAND2X1 U748 ( .A(n1029), .B(n2018), .Y(n1027) );
  ADDFX1 U749 ( .A(n1299), .B(n1300), .CI(n1298), .CO(n1350), .S(n1305) );
  OAI2BB1X2 U750 ( .A0N(n1109), .A1N(n3364), .B0(n1108), .Y(n3358) );
  ADDFX1 U751 ( .A(n3020), .B(n3019), .CI(n3018), .CO(n3049), .S(n3163) );
  ADDFX2 U752 ( .A(n1373), .B(n1372), .CI(n1371), .CO(n1382), .S(n1399) );
  ADDFX1 U753 ( .A(n2721), .B(n2720), .CI(n2719), .CO(n3438), .S(n2709) );
  ADDFX1 U754 ( .A(n1309), .B(n1308), .CI(n1307), .CO(n1306), .S(n1386) );
  ADDFX1 U755 ( .A(n1403), .B(n1402), .CI(n1401), .CO(n1441), .S(n1445) );
  ADDFX1 U756 ( .A(n3318), .B(n3317), .CI(n3316), .CO(n3319), .S(n3309) );
  ADDFHX1 U757 ( .A(n3083), .B(n3081), .CI(n3082), .CO(n3126), .S(n3099) );
  ADDFHX1 U758 ( .A(n3233), .B(n3232), .CI(n3231), .CO(n3226), .S(n3315) );
  ADDFX1 U759 ( .A(n2546), .B(n2545), .CI(n2544), .CO(n2658), .S(n2521) );
  OAI2BB1X1 U760 ( .A0N(n2548), .A1N(n1104), .B0(n1103), .Y(n2523) );
  ADDFX2 U761 ( .A(n2919), .B(n2920), .CI(n2921), .CO(n3342), .S(n3361) );
  OAI2BB1X1 U762 ( .A0N(n766), .A1N(n2916), .B0(n765), .Y(n3340) );
  ADDFX1 U763 ( .A(n2256), .B(n2255), .CI(n2254), .CO(n2311), .S(n2252) );
  ADDFX1 U764 ( .A(n3221), .B(n3220), .CI(n3219), .CO(n3222), .S(n3241) );
  ADDFX1 U765 ( .A(n3214), .B(n3176), .CI(n3213), .CO(n3223), .S(n3243) );
  OAI22X1 U766 ( .A0(n3053), .A1(n3259), .B0(n3052), .B1(n3261), .Y(n3083) );
  OAI2BB1X1 U767 ( .A0N(n817), .A1N(n2108), .B0(n816), .Y(n2159) );
  NAND2X1 U768 ( .A(n1938), .B(n1937), .Y(n2042) );
  OAI2BB2X2 U769 ( .B0(n3067), .B1(n3179), .A0N(n677), .A1N(n676), .Y(n3081)
         );
  ADDFHX1 U770 ( .A(n1808), .B(n1807), .CI(n1806), .CO(n1822), .S(n1843) );
  ADDFHX1 U771 ( .A(n1512), .B(n1511), .CI(n1510), .CO(n1553), .S(n1501) );
  XNOR2X1 U772 ( .A(n3173), .B(n3054), .Y(n3067) );
  ADDHXL U773 ( .A(n2992), .B(n2991), .CO(n3025), .S(n3198) );
  OR2XL U774 ( .A(n2789), .B(n3110), .Y(n1098) );
  OAI22X1 U775 ( .A0(n3069), .A1(n3070), .B0(n3056), .B1(n3068), .Y(n3101) );
  NAND2X1 U776 ( .A(n860), .B(n857), .Y(n3034) );
  ADDFHX1 U777 ( .A(n2559), .B(n2558), .CI(n2557), .CO(n2552), .S(n2597) );
  ADDFHX1 U778 ( .A(n3074), .B(n3073), .CI(n3072), .CO(n3123), .S(n3134) );
  ADDFX1 U779 ( .A(n2538), .B(n2537), .CI(n2536), .CO(n2655), .S(n2533) );
  BUFX2 U780 ( .A(n3451), .Y(n755) );
  ADDHXL U781 ( .A(n1076), .B(n1538), .CO(n1584), .S(n1561) );
  OR2XL U782 ( .A(n2781), .B(n2782), .Y(n2775) );
  XNOR2XL U783 ( .A(n1038), .B(n1791), .Y(n1324) );
  OR2X1 U784 ( .A(n2482), .B(n2481), .Y(n2542) );
  AND2X1 U785 ( .A(n2630), .B(n2629), .Y(n1050) );
  OR2X1 U786 ( .A(n2163), .B(n2162), .Y(n2217) );
  XOR2X1 U787 ( .A(n3251), .B(n587), .Y(n1287) );
  OR2XL U788 ( .A(n2968), .B(n3182), .Y(n860) );
  OR2X1 U789 ( .A(n1888), .B(n1887), .Y(n1933) );
  ADDFX2 U790 ( .A(n3282), .B(n3281), .CI(n3280), .CO(n3305), .S(n3288) );
  OAI2BB2X1 U791 ( .B0(n2934), .B1(n3087), .A0N(n732), .A1N(n3084), .Y(n3074)
         );
  OAI2BB2X1 U792 ( .B0(n1540), .B1(n1607), .A0N(n634), .A1N(n1606), .Y(n1583)
         );
  OAI22X1 U793 ( .A0(n2931), .A1(n3068), .B0(n2882), .B1(n3070), .Y(n2917) );
  ADDFHX1 U794 ( .A(n2813), .B(n2812), .CI(n2811), .CO(n2809), .S(n2822) );
  ADDFX2 U795 ( .A(n2239), .B(n2238), .CI(n2237), .CO(n2253), .S(n2235) );
  OAI2BB1XL U796 ( .A0N(n683), .A1N(n1009), .B0(n1008), .Y(n2813) );
  BUFX4 U797 ( .A(n3004), .Y(n1017) );
  ADDFX1 U798 ( .A(n2804), .B(n2803), .CI(n2802), .CO(n2819), .S(n2814) );
  BUFX4 U799 ( .A(n972), .Y(n773) );
  OAI22X1 U800 ( .A0(n1776), .A1(n2264), .B0(n2263), .B1(n697), .Y(n1801) );
  ADDFHX1 U801 ( .A(n2516), .B(n2517), .CI(n2515), .CO(n2549), .S(n2585) );
  ADDFHX1 U802 ( .A(n2520), .B(n2519), .CI(n2518), .CO(n2548), .S(n2584) );
  AND2X1 U803 ( .A(n645), .B(n2971), .Y(n2973) );
  NAND2BX2 U804 ( .AN(n3270), .B(n1954), .Y(n1333) );
  INVX2 U805 ( .A(n1954), .Y(n573) );
  INVX2 U806 ( .A(n3237), .Y(n590) );
  XNOR2X1 U807 ( .A(n2888), .B(n1242), .Y(n1243) );
  BUFX4 U808 ( .A(n1235), .Y(n3179) );
  OAI22X1 U809 ( .A0(n2458), .A1(n4082), .B0(n2429), .B1(n4081), .Y(n2519) );
  OAI22X1 U810 ( .A0(n2913), .A1(n3182), .B0(n2835), .B1(n3184), .Y(n2903) );
  NOR2BX1 U811 ( .AN(n3270), .B(n3446), .Y(n2615) );
  BUFX12 U812 ( .A(n2569), .Y(n3239) );
  BUFX2 U813 ( .A(n1202), .Y(n1606) );
  OR2XL U814 ( .A(n2006), .B(n2126), .Y(n636) );
  OR2XL U815 ( .A(n2618), .B(n2755), .Y(n896) );
  NAND2X1 U816 ( .A(n1062), .B(n1060), .Y(n1059) );
  NAND2X2 U817 ( .A(n2974), .B(n3275), .Y(n3273) );
  XOR2X2 U818 ( .A(n2890), .B(n2889), .Y(n3261) );
  BUFX8 U819 ( .A(n3166), .Y(n769) );
  XOR2X1 U820 ( .A(n2975), .B(n2900), .Y(n1062) );
  XOR2X2 U821 ( .A(n3251), .B(n2197), .Y(n815) );
  NAND2X2 U822 ( .A(n1701), .B(n1183), .Y(n1700) );
  BUFX2 U823 ( .A(n3237), .Y(n3253) );
  NOR2X1 U824 ( .A(n2892), .B(butt_a_real[1]), .Y(n2884) );
  XNOR2X1 U825 ( .A(n2506), .B(n2499), .Y(n2503) );
  BUFX16 U826 ( .A(n2783), .Y(n3251) );
  XNOR2X1 U827 ( .A(butt_b_imag[4]), .B(butt_a_imag[4]), .Y(n1226) );
  XNOR2X1 U828 ( .A(n2425), .B(n2418), .Y(n2422) );
  XNOR2X1 U829 ( .A(n2746), .B(n2739), .Y(n2743) );
  NAND2X2 U830 ( .A(n2199), .B(n1637), .Y(n2198) );
  NAND2X2 U831 ( .A(n1200), .B(n717), .Y(n2788) );
  NAND2X2 U832 ( .A(n1068), .B(n2639), .Y(n2502) );
  XNOR3X2 U833 ( .A(n1191), .B(n2632), .C(n952), .Y(n1793) );
  XNOR2XL U834 ( .A(n2453), .B(n1787), .Y(n1790) );
  XNOR2X2 U835 ( .A(n2462), .B(n2461), .Y(n2432) );
  XNOR2X2 U836 ( .A(n2455), .B(n1951), .Y(n1880) );
  INVX4 U837 ( .A(n805), .Y(n3112) );
  XOR2X2 U838 ( .A(n2750), .B(n1018), .Y(n3181) );
  NAND2X1 U839 ( .A(n1575), .B(n1574), .Y(n1576) );
  XNOR2X1 U840 ( .A(n1520), .B(n1474), .Y(n1478) );
  XOR2X1 U841 ( .A(n1656), .B(butt_a_imag[12]), .Y(n1658) );
  XOR2X1 U842 ( .A(n1069), .B(n2639), .Y(n3028) );
  OAI21X2 U843 ( .A0(butt_b_imag[10]), .A1(n1035), .B0(n1034), .Y(n1574) );
  OAI2BB1X1 U844 ( .A0N(butt_a_real[4]), .A1N(n2744), .B0(n2633), .Y(n2750) );
  XOR2X1 U845 ( .A(n1518), .B(butt_a_imag[10]), .Y(n1520) );
  OAI21X2 U846 ( .A0(n1089), .A1(n1088), .B0(n1150), .Y(n1220) );
  NAND2X1 U847 ( .A(n1272), .B(n1271), .Y(n997) );
  XOR2X1 U848 ( .A(butt_b_imag[11]), .B(butt_a_imag[11]), .Y(n1575) );
  NAND2X1 U849 ( .A(n915), .B(n832), .Y(n831) );
  NAND2XL U850 ( .A(n1224), .B(butt_a_imag[4]), .Y(n1150) );
  BUFX8 U851 ( .A(n1193), .Y(n1261) );
  XOR2X1 U852 ( .A(n1892), .B(butt_a_imag[16]), .Y(n1894) );
  XNOR2X1 U853 ( .A(n1166), .B(n2057), .Y(n1249) );
  BUFX2 U854 ( .A(n1167), .Y(n1168) );
  INVX2 U855 ( .A(n1140), .Y(n925) );
  INVX2 U856 ( .A(lay_cnt[5]), .Y(n4640) );
  NAND2X1 U857 ( .A(n2072), .B(lay_cnt[4]), .Y(n1137) );
  INVX2 U858 ( .A(n3817), .Y(n678) );
  NOR2X1 U859 ( .A(n3812), .B(n3840), .Y(n1135) );
  INVXL U860 ( .A(butt_b_real[14]), .Y(n2465) );
  BUFX1 U861 ( .A(n2453), .Y(n733) );
  INVXL U862 ( .A(n2711), .Y(n574) );
  INVXL U863 ( .A(n3028), .Y(n973) );
  XOR2XL U864 ( .A(n645), .B(n3028), .Y(n2985) );
  INVXL U865 ( .A(n1476), .Y(n808) );
  XOR2XL U866 ( .A(n2897), .B(n2894), .Y(n2895) );
  NOR2XL U867 ( .A(n2009), .B(butt_a_imag[17]), .Y(n922) );
  XNOR2XL U868 ( .A(n580), .B(n657), .Y(n2026) );
  XNOR2XL U869 ( .A(n3234), .B(n657), .Y(n1973) );
  XNOR2XL U870 ( .A(n3250), .B(n657), .Y(n1799) );
  NAND2X1 U871 ( .A(n951), .B(n1791), .Y(n1887) );
  NAND2X1 U872 ( .A(n878), .B(n877), .Y(n876) );
  INVXL U873 ( .A(n2413), .Y(n2674) );
  XNOR2XL U874 ( .A(n2976), .B(n2567), .Y(n2698) );
  XNOR2XL U875 ( .A(n645), .B(n2757), .Y(n2758) );
  XNOR2XL U876 ( .A(n3009), .B(n3181), .Y(n3089) );
  XNOR2XL U877 ( .A(n2976), .B(n594), .Y(n2987) );
  XNOR2XL U878 ( .A(n3054), .B(n3253), .Y(n3011) );
  XNOR2XL U879 ( .A(n3014), .B(n2979), .Y(n1591) );
  XOR3X2 U880 ( .A(n1000), .B(n1338), .C(n997), .Y(n805) );
  INVXL U881 ( .A(n3258), .Y(n588) );
  XOR2XL U882 ( .A(n1073), .B(n590), .Y(n3168) );
  OAI22X1 U883 ( .A0(n2969), .A1(n3112), .B0(n3110), .B1(n1041), .Y(n996) );
  INVXL U884 ( .A(butt_b_real[17]), .Y(n2409) );
  XNOR2XL U885 ( .A(n3054), .B(n1749), .Y(n2181) );
  AOI2BB1X1 U886 ( .A0N(n2205), .A1N(n3558), .B0(n828), .Y(n827) );
  NAND2X1 U887 ( .A(n636), .B(n637), .Y(n2112) );
  XNOR2XL U888 ( .A(n745), .B(n1606), .Y(n1408) );
  ADDHX1 U889 ( .A(n1801), .B(n1800), .CO(n1916), .S(n1831) );
  XNOR2XL U890 ( .A(n2976), .B(n4076), .Y(n3441) );
  XNOR2XL U891 ( .A(n1643), .B(n1642), .Y(n1682) );
  ADDFX2 U892 ( .A(n2562), .B(n2561), .CI(n2560), .CO(n2582), .S(n2596) );
  NOR2XL U893 ( .A(n4275), .B(n4277), .Y(n3476) );
  XNOR2XL U894 ( .A(n2976), .B(n1173), .Y(n1592) );
  XNOR2XL U895 ( .A(n580), .B(n3173), .Y(n1326) );
  NAND2X1 U896 ( .A(n1252), .B(n3271), .Y(n3269) );
  XOR2XL U897 ( .A(n3488), .B(n2001), .Y(n2002) );
  ADDFX2 U898 ( .A(n2038), .B(n2037), .CI(n2036), .CO(n2137), .S(n2035) );
  NOR2XL U899 ( .A(n3736), .B(n3731), .Y(n3725) );
  ADDFX2 U900 ( .A(n3171), .B(n3170), .CI(n3169), .CO(n3161), .S(n3207) );
  NOR2XL U901 ( .A(Q[7]), .B(butt_a_imag[7]), .Y(n4054) );
  XOR2X1 U902 ( .A(n2193), .B(n2194), .Y(n2186) );
  NOR2XL U903 ( .A(Q[32]), .B(butt_a_real[13]), .Y(n3982) );
  NAND2X1 U904 ( .A(n3422), .B(n3421), .Y(n3474) );
  NOR2XL U905 ( .A(Q[25]), .B(butt_a_real[6]), .Y(n4335) );
  ADDFHX1 U906 ( .A(n3127), .B(n3126), .CI(n3125), .CO(n3368), .S(n3152) );
  INVXL U907 ( .A(n3542), .Y(n3556) );
  NOR2XL U908 ( .A(Q[6]), .B(butt_a_imag[6]), .Y(n4052) );
  NOR2XL U909 ( .A(Q[34]), .B(butt_a_real[15]), .Y(n4446) );
  ADDFXL U910 ( .A(n4653), .B(n4673), .CI(n4089), .CO(n4090), .S(n4527) );
  OR2X2 U911 ( .A(n1468), .B(n1469), .Y(n3680) );
  NOR2X2 U912 ( .A(n647), .B(n4035), .Y(n4042) );
  AND2X1 U913 ( .A(n3690), .B(n3689), .Y(n3691) );
  XOR2X1 U914 ( .A(n833), .B(n1117), .Y(n3581) );
  XNOR2X1 U915 ( .A(n2327), .B(n2326), .Y(n4214) );
  INVXL U916 ( .A(n4184), .Y(n4186) );
  XNOR2XL U917 ( .A(n3904), .B(n3903), .Y(n4359) );
  INVXL U918 ( .A(Q[11]), .Y(n3885) );
  INVXL U919 ( .A(Q[23]), .Y(n3863) );
  INVXL U920 ( .A(Q[34]), .Y(n3884) );
  NOR2XL U921 ( .A(n4102), .B(lay_cnt[0]), .Y(N1236) );
  INVXL U922 ( .A(n1046), .Y(n596) );
  AND2X2 U923 ( .A(n4652), .B(n3859), .Y(n570) );
  INVXL U924 ( .A(n4145), .Y(n4147) );
  NOR2X1 U925 ( .A(n4677), .B(lay_cnt[1]), .Y(n4145) );
  BUFX2 U926 ( .A(n1190), .Y(n1791) );
  INVX2 U927 ( .A(n2821), .Y(n1095) );
  INVXL U928 ( .A(n735), .Y(n1030) );
  XOR3X2 U929 ( .A(n3370), .B(n3372), .C(n3371), .Y(n3405) );
  NAND2X1 U930 ( .A(n880), .B(n3410), .Y(n3600) );
  INVXL U931 ( .A(n710), .Y(n3629) );
  BUFX2 U932 ( .A(n1252), .Y(n594) );
  INVX2 U933 ( .A(n1079), .Y(n3256) );
  NAND2X1 U934 ( .A(n3581), .B(n4598), .Y(n3587) );
  NAND4X1 U935 ( .A(n4205), .B(n4204), .C(n4203), .D(n4202), .Y(D_imag[12]) );
  NAND4X1 U936 ( .A(n4445), .B(n4444), .C(n4443), .D(n4442), .Y(D_real[11]) );
  NAND4X1 U937 ( .A(n3993), .B(n3994), .C(n3995), .D(n3992), .Y(D_real[12]) );
  NAND2XL U938 ( .A(n4214), .B(n4594), .Y(n2334) );
  OAI211X1 U939 ( .A0(n4593), .A1(n4592), .B0(n4590), .C0(n4591), .Y(D_imag[7]) );
  NAND2XL U940 ( .A(n4214), .B(n4598), .Y(n4217) );
  NAND2XL U941 ( .A(n4433), .B(n4614), .Y(n746) );
  AOI21XL U942 ( .A0(n4598), .A1(n4572), .B0(n3685), .Y(n3686) );
  OAI2BB1X1 U943 ( .A0N(n4594), .A1N(n4573), .B0(n4261), .Y(D_imag[1]) );
  OAI211X1 U944 ( .A0(n3930), .A1(n4270), .B0(n3929), .C0(n3928), .Y(D_real[0]) );
  CLKBUFX1 U945 ( .A(n3967), .Y(n3969) );
  INVX1 U946 ( .A(n4308), .Y(n4321) );
  NOR2X1 U947 ( .A(n820), .B(n2338), .Y(n2322) );
  AOI21X1 U948 ( .A0(n2374), .A1(n2278), .B0(n2373), .Y(n2375) );
  OAI211X1 U949 ( .A0(n3962), .A1(n4270), .B0(n3961), .C0(n3960), .Y(D_imag[0]) );
  INVX1 U950 ( .A(n3997), .Y(n4028) );
  INVX1 U951 ( .A(n2146), .Y(n2374) );
  INVX1 U952 ( .A(n2343), .Y(n2325) );
  AOI21X1 U953 ( .A0(n2343), .A1(n2342), .B0(n2341), .Y(n964) );
  BUFXL U954 ( .A(n3650), .Y(n4032) );
  ADDFHX2 U955 ( .A(n2145), .B(n2144), .CI(n2143), .CO(n2275), .S(n2052) );
  INVX3 U956 ( .A(n3473), .Y(n571) );
  NOR2X2 U957 ( .A(n880), .B(n3410), .Y(n4324) );
  NAND2X2 U958 ( .A(n3404), .B(n3403), .Y(n3592) );
  AND2X1 U959 ( .A(n3469), .B(n3468), .Y(n1120) );
  BUFXL U960 ( .A(n3902), .Y(n650) );
  NAND2BX2 U961 ( .AN(n3429), .B(n702), .Y(n3469) );
  NAND2X2 U962 ( .A(n1865), .B(n1864), .Y(n3640) );
  ADDFHX2 U963 ( .A(n1860), .B(n1859), .CI(n1858), .CO(n1871), .S(n1868) );
  INVX2 U964 ( .A(n3583), .Y(n3548) );
  NAND2X2 U965 ( .A(n3630), .B(n4310), .Y(n958) );
  INVX1 U966 ( .A(n3332), .Y(n855) );
  NAND2X1 U967 ( .A(n2370), .B(n2369), .Y(n3582) );
  ADDFHX2 U968 ( .A(n2727), .B(n2726), .CI(n2725), .CO(n3425), .S(n3423) );
  INVX1 U969 ( .A(n3508), .Y(n4068) );
  AND2XL U970 ( .A(n4088), .B(n4508), .Y(n1113) );
  NAND2XL U971 ( .A(n918), .B(n735), .Y(n1028) );
  NAND2XL U972 ( .A(n2249), .B(n2250), .Y(n758) );
  INVX1 U973 ( .A(n3547), .Y(n3585) );
  NAND2X1 U974 ( .A(n3457), .B(n3456), .Y(n4069) );
  NAND2X1 U975 ( .A(n3327), .B(n3326), .Y(n4309) );
  INVX1 U976 ( .A(n1027), .Y(n918) );
  NAND2XL U977 ( .A(n2810), .B(n1048), .Y(n1047) );
  INVX3 U978 ( .A(n638), .Y(n639) );
  AND2XL U979 ( .A(n4521), .B(n4520), .Y(n1119) );
  INVXL U980 ( .A(n2822), .Y(n625) );
  ADDFHX2 U981 ( .A(n2236), .B(n2235), .CI(n2234), .CO(n2272), .S(n2248) );
  ADDFHX2 U982 ( .A(n2724), .B(n2723), .CI(n2722), .CO(n3435), .S(n2706) );
  NAND2X1 U983 ( .A(n705), .B(n1042), .Y(n2869) );
  OAI21XL U984 ( .A0(n3034), .A1(n3035), .B0(n3033), .Y(n3037) );
  ADDFHX2 U985 ( .A(n1616), .B(n1615), .CI(n1614), .CO(n1736), .S(n1598) );
  ADDFX1 U986 ( .A(n4075), .B(n4074), .CI(n4073), .CO(n4087), .S(n3522) );
  OAI2BB1X2 U987 ( .A0N(n1092), .A1N(n1487), .B0(n1091), .Y(n1537) );
  ADDFHX2 U988 ( .A(n2221), .B(n2220), .CI(n2219), .CO(n2225), .S(n2191) );
  ADDFX1 U989 ( .A(n3298), .B(n3297), .CI(n3296), .CO(n3318), .S(n3291) );
  AND2XL U990 ( .A(n1427), .B(n1426), .Y(n1428) );
  AND2XL U991 ( .A(n1418), .B(n1417), .Y(n1419) );
  NAND2XL U992 ( .A(n3022), .B(n686), .Y(n685) );
  ADDFHX1 U993 ( .A(n1306), .B(n1305), .CI(n1304), .CO(n1347), .S(n1370) );
  NAND2XL U994 ( .A(n991), .B(n989), .Y(n3146) );
  ADDFHX2 U995 ( .A(n2853), .B(n2852), .CI(n2851), .CO(n2823), .S(n3338) );
  CLKINVX2 U996 ( .A(n2824), .Y(n1043) );
  AND2XL U997 ( .A(n3278), .B(n3277), .Y(n3279) );
  OR2XL U998 ( .A(n2928), .B(n3112), .Y(n991) );
  NAND2XL U999 ( .A(n2549), .B(n2550), .Y(n1103) );
  ADDFHX1 U1000 ( .A(n3080), .B(n3079), .CI(n3078), .CO(n3122), .S(n3127) );
  XOR2X2 U1001 ( .A(n1010), .B(n1009), .Y(n2794) );
  NAND2X1 U1002 ( .A(n2990), .B(n2989), .Y(n1022) );
  CLKBUFX1 U1003 ( .A(n1684), .Y(n656) );
  INVX2 U1004 ( .A(n876), .Y(n874) );
  ADDFHX2 U1005 ( .A(n1877), .B(n1876), .CI(n1875), .CO(n1979), .S(n1919) );
  NAND2X2 U1006 ( .A(n797), .B(n794), .Y(n1345) );
  OAI22X1 U1007 ( .A0(n2970), .A1(n3070), .B0(n975), .B1(n3068), .Y(n3039) );
  OR2X2 U1008 ( .A(n1778), .B(n2198), .Y(n849) );
  OR2XL U1009 ( .A(n2554), .B(n2555), .Y(n2515) );
  NAND2BXL U1010 ( .AN(n3239), .B(n2830), .Y(n1671) );
  NAND2BXL U1011 ( .AN(n3239), .B(n2979), .Y(n1241) );
  NAND2BXL U1012 ( .AN(n645), .B(n2674), .Y(n2414) );
  BUFX12 U1013 ( .A(n2788), .Y(n3054) );
  BUFX12 U1014 ( .A(n2733), .Y(n3164) );
  NAND2X1 U1015 ( .A(n887), .B(n1216), .Y(n1217) );
  AOI21XL U1016 ( .A0(n3493), .A1(n3491), .B0(n3486), .Y(n3487) );
  OAI2BB1X1 U1017 ( .A0N(n4623), .A1N(n4627), .B0(n4649), .Y(n3856) );
  INVX2 U1018 ( .A(n4563), .Y(n4605) );
  NAND2X1 U1019 ( .A(n915), .B(n888), .Y(n887) );
  INVXL U1020 ( .A(n3444), .Y(n2721) );
  INVX3 U1021 ( .A(n915), .Y(n830) );
  INVX2 U1022 ( .A(n4594), .Y(n4592) );
  INVX2 U1023 ( .A(n4661), .Y(n4664) );
  INVX2 U1024 ( .A(n2071), .Y(n4552) );
  INVX1 U1025 ( .A(n3821), .Y(n4106) );
  NAND2X1 U1026 ( .A(n3799), .B(n3806), .Y(n3768) );
  INVXL U1027 ( .A(n1955), .Y(n611) );
  NOR2X4 U1028 ( .A(n2371), .B(n4502), .Y(n4598) );
  NOR2X4 U1029 ( .A(n2371), .B(n2332), .Y(n4596) );
  INVXL U1030 ( .A(n592), .Y(n615) );
  CLKBUFX1 U1031 ( .A(n2055), .Y(n3798) );
  INVX2 U1032 ( .A(n591), .Y(n572) );
  NAND2X1 U1033 ( .A(in_out_cnt[6]), .B(n4659), .Y(n4657) );
  INVX2 U1034 ( .A(n657), .Y(n592) );
  OAI2BB1XL U1035 ( .A0N(butt_b_real[8]), .A1N(n4186), .B0(n4158), .Y(n520) );
  NAND2BXL U1036 ( .AN(n1339), .B(n810), .Y(n809) );
  NAND2XL U1037 ( .A(n2435), .B(n1604), .Y(n1605) );
  NAND2X1 U1038 ( .A(IN_VALID), .B(n2081), .Y(n4669) );
  INVX2 U1039 ( .A(n594), .Y(n575) );
  INVX2 U1040 ( .A(n3028), .Y(n576) );
  NAND2BXL U1041 ( .AN(n1250), .B(n1249), .Y(n1083) );
  INVX2 U1042 ( .A(n3866), .Y(n653) );
  NAND2BXL U1043 ( .AN(n1197), .B(n979), .Y(n955) );
  NAND2X1 U1044 ( .A(n2403), .B(n2402), .Y(n2413) );
  NAND2X1 U1045 ( .A(in_out_cnt[4]), .B(n4656), .Y(n4654) );
  NAND2X1 U1046 ( .A(n1648), .B(n1647), .Y(n1655) );
  XNOR2X1 U1047 ( .A(n2467), .B(n2460), .Y(n2464) );
  INVX2 U1048 ( .A(n1272), .Y(n1031) );
  OAI21XL U1049 ( .A0(n2634), .A1(butt_a_real[6]), .B0(butt_a_real[5]), .Y(
        n2501) );
  INVX2 U1050 ( .A(n2751), .Y(n1018) );
  INVXL U1051 ( .A(n3891), .Y(n629) );
  NAND2XL U1052 ( .A(n2465), .B(butt_a_real[14]), .Y(n2447) );
  INVXL U1053 ( .A(n3860), .Y(n632) );
  INVXL U1054 ( .A(n3877), .Y(n633) );
  NAND2XL U1055 ( .A(n1766), .B(butt_a_imag[14]), .Y(n1759) );
  INVX2 U1056 ( .A(mode_val), .Y(n3858) );
  INVX2 U1057 ( .A(Q[21]), .Y(n3896) );
  INVX2 U1058 ( .A(Q[22]), .Y(n3892) );
  INVX2 U1059 ( .A(Q[20]), .Y(n3894) );
  INVX2 U1060 ( .A(Q[3]), .Y(n3891) );
  INVX2 U1061 ( .A(Q[19]), .Y(n3868) );
  INVX2 U1062 ( .A(Q[24]), .Y(n3870) );
  INVX2 U1063 ( .A(Q[25]), .Y(n3872) );
  INVX2 U1064 ( .A(Q[36]), .Y(n3888) );
  NAND2X1 U1065 ( .A(rst_n), .B(OUT_VALID), .Y(n3857) );
  INVX2 U1066 ( .A(Q[26]), .Y(n3874) );
  INVX2 U1067 ( .A(Q[18]), .Y(n4652) );
  INVX2 U1068 ( .A(Q[8]), .Y(n3860) );
  INVX2 U1069 ( .A(Q[35]), .Y(n3876) );
  INVX2 U1070 ( .A(butt_b_real[12]), .Y(n2436) );
  INVX2 U1071 ( .A(Q[27]), .Y(n3861) );
  INVX2 U1072 ( .A(Q[9]), .Y(n3877) );
  INVX2 U1073 ( .A(Q[28]), .Y(n3878) );
  INVX2 U1074 ( .A(butt_b_imag[1]), .Y(n1166) );
  INVX2 U1075 ( .A(Q[33]), .Y(n3882) );
  INVX2 U1076 ( .A(Q[10]), .Y(n3889) );
  INVX2 U1077 ( .A(Q[32]), .Y(n3880) );
  INVX2 U1078 ( .A(Q[29]), .Y(n3890) );
  INVX2 U1079 ( .A(Q[30]), .Y(n3886) );
  INVX2 U1080 ( .A(Q[31]), .Y(n3865) );
  INVX1 U1081 ( .A(Q[4]), .Y(n3862) );
  INVX1 U1082 ( .A(Q[5]), .Y(n3869) );
  INVX1 U1083 ( .A(Q[6]), .Y(n3871) );
  XNOR2X2 U1084 ( .A(butt_a_real[6]), .B(butt_b_real[6]), .Y(n2632) );
  INVX1 U1085 ( .A(Q[7]), .Y(n3873) );
  INVX1 U1086 ( .A(Q[1]), .Y(n3893) );
  INVX2 U1087 ( .A(butt_a_imag[3]), .Y(n1088) );
  XNOR2X2 U1088 ( .A(butt_b_real[8]), .B(butt_a_real[8]), .Y(n2506) );
  INVX1 U1089 ( .A(Q[12]), .Y(n3864) );
  INVX1 U1090 ( .A(Q[13]), .Y(n3879) );
  CLKBUFX1 U1091 ( .A(Q[14]), .Y(n3881) );
  CLKBUFX1 U1092 ( .A(Q[17]), .Y(n3887) );
  INVX2 U1093 ( .A(is_row), .Y(n4644) );
  CLKBUFX1 U1094 ( .A(Q[15]), .Y(n3883) );
  NAND2X1 U1095 ( .A(n4504), .B(n4598), .Y(n3524) );
  NAND2X1 U1096 ( .A(n621), .B(n1119), .Y(n624) );
  INVX1 U1097 ( .A(n889), .Y(n600) );
  XNOR2X2 U1098 ( .A(n2319), .B(n2318), .Y(n4230) );
  XOR2X2 U1099 ( .A(n791), .B(n663), .Y(n4504) );
  NAND2X1 U1100 ( .A(n4097), .B(n3459), .Y(n4503) );
  XOR2X2 U1101 ( .A(n3973), .B(n1116), .Y(n4532) );
  XNOR2X2 U1102 ( .A(n4474), .B(n4473), .Y(n4490) );
  NAND2XL U1103 ( .A(n655), .B(n4594), .Y(n4065) );
  OAI2BB1X1 U1104 ( .A0N(n4594), .A1N(n4615), .B0(n3686), .Y(D_imag[4]) );
  OAI2BB1X1 U1105 ( .A0N(n4594), .A1N(n4359), .B0(n4290), .Y(D_real[1]) );
  OAI2BB1X1 U1106 ( .A0N(n4598), .A1N(n4308), .B0(n4307), .Y(D_real[2]) );
  XOR2X2 U1107 ( .A(n737), .B(n662), .Y(n4599) );
  XOR2X2 U1108 ( .A(n4383), .B(n1121), .Y(n879) );
  NOR2X1 U1109 ( .A(n1123), .B(n4541), .Y(n4317) );
  XOR2X2 U1110 ( .A(n692), .B(n3691), .Y(n4597) );
  XOR2X1 U1111 ( .A(n3603), .B(n3602), .Y(n4410) );
  NOR2X1 U1112 ( .A(n1123), .B(n4270), .Y(n4289) );
  XOR2X1 U1113 ( .A(n4333), .B(n4332), .Y(n4441) );
  OAI2BB1X1 U1114 ( .A0N(n4598), .A1N(n4432), .B0(n4431), .Y(D_imag[2]) );
  INVX1 U1115 ( .A(n4432), .Y(n4551) );
  XOR2X1 U1116 ( .A(n3653), .B(n3652), .Y(n4572) );
  NOR2X1 U1117 ( .A(n4587), .B(n4541), .Y(n4547) );
  NOR2X1 U1118 ( .A(n4587), .B(n4270), .Y(n4260) );
  NOR2X1 U1119 ( .A(n4587), .B(n4592), .Y(n4430) );
  OAI21X2 U1120 ( .A0(n2344), .A1(n2345), .B0(n964), .Y(n1053) );
  INVX1 U1121 ( .A(n3898), .Y(n4264) );
  NOR2X1 U1122 ( .A(n4322), .B(n721), .Y(n4328) );
  INVX4 U1123 ( .A(n3976), .Y(n577) );
  INVXL U1124 ( .A(n4511), .Y(n4512) );
  ADDFHX2 U1125 ( .A(n2224), .B(n2223), .CI(n2222), .CO(n2284), .S(n2282) );
  NOR2X1 U1126 ( .A(n4506), .B(n4509), .Y(n4507) );
  XNOR3X2 U1127 ( .A(n1857), .B(n1856), .C(n1855), .Y(n1858) );
  AOI2BB1X2 U1128 ( .A0N(n3330), .A1N(n4309), .B0(n3629), .Y(n957) );
  INVX3 U1129 ( .A(n3957), .Y(n939) );
  OAI2BB1X2 U1130 ( .A0N(n1924), .A1N(n841), .B0(n839), .Y(n1965) );
  NAND2X2 U1131 ( .A(n1624), .B(n1623), .Y(n3957) );
  OAI2BB1X2 U1132 ( .A0N(n1028), .A1N(n2138), .B0(n1026), .Y(n2156) );
  NOR2X1 U1133 ( .A(n2370), .B(n2369), .Y(n3583) );
  INVX2 U1134 ( .A(n2154), .Y(n2139) );
  ADDFHX2 U1135 ( .A(n2730), .B(n2729), .CI(n2728), .CO(n3428), .S(n3426) );
  ADDFHX2 U1136 ( .A(n1928), .B(n1927), .CI(n1926), .CO(n1983), .S(n1929) );
  ADDFHX2 U1137 ( .A(n2707), .B(n2706), .CI(n2705), .CO(n3430), .S(n3427) );
  CLKINVX2 U1138 ( .A(n3209), .Y(n4310) );
  OAI2BB1X2 U1139 ( .A0N(n1049), .A1N(n2809), .B0(n1047), .Y(n2956) );
  NOR2X1 U1140 ( .A(n3329), .B(n3328), .Y(n3330) );
  AND2X1 U1141 ( .A(n3566), .B(n3569), .Y(n1112) );
  NAND2X1 U1142 ( .A(n1467), .B(n1466), .Y(n4537) );
  XNOR3X2 U1143 ( .A(n1925), .B(n1924), .C(n843), .Y(n1931) );
  NOR2X1 U1144 ( .A(n3457), .B(n3456), .Y(n3508) );
  ADDFHX2 U1145 ( .A(n3121), .B(n3119), .CI(n3120), .CO(n3334), .S(n3331) );
  ADDFHX2 U1146 ( .A(n2137), .B(n2136), .CI(n2135), .CO(n2154), .S(n2141) );
  ADDFHX2 U1147 ( .A(n2296), .B(n2295), .CI(n2294), .CO(n2317), .S(n2286) );
  NAND2BXL U1148 ( .AN(n3159), .B(n709), .Y(n708) );
  ADDFHX2 U1149 ( .A(n1982), .B(n1981), .CI(n1980), .CO(n2030), .S(n1985) );
  ADDFHX2 U1150 ( .A(n2192), .B(n2191), .CI(n2190), .CO(n2224), .S(n2196) );
  ADDFHX2 U1151 ( .A(n3139), .B(n3138), .CI(n3137), .CO(n3401), .S(n3155) );
  NAND2X1 U1152 ( .A(n626), .B(n2820), .Y(n960) );
  ADDFHX2 U1153 ( .A(n2523), .B(n2522), .CI(n2521), .CO(n2727), .S(n2601) );
  ADDFHX2 U1154 ( .A(n2650), .B(n2649), .CI(n2648), .CO(n2654), .S(n2958) );
  ADDFHX2 U1155 ( .A(n2273), .B(n2272), .CI(n2271), .CO(n2294), .S(n2249) );
  NOR2X1 U1156 ( .A(n3550), .B(n3549), .Y(n3547) );
  ADDFHX2 U1157 ( .A(n1370), .B(n1369), .CI(n1368), .CO(n1466), .S(n1462) );
  ADDFHX2 U1158 ( .A(n1619), .B(n1618), .CI(n1617), .CO(n1735), .S(n1622) );
  NAND2X2 U1159 ( .A(n907), .B(n906), .Y(n2703) );
  ADDFHX2 U1160 ( .A(n3192), .B(n3191), .CI(n3190), .CO(n3328), .S(n3327) );
  ADDFHX2 U1161 ( .A(n1366), .B(n1367), .CI(n1365), .CO(n1469), .S(n1467) );
  ADDFHX2 U1162 ( .A(n2682), .B(n2681), .CI(n2680), .CO(n2728), .S(n2725) );
  ADDFHX2 U1163 ( .A(n1568), .B(n1569), .CI(n1567), .CO(n1597), .S(n1572) );
  ADDFHX2 U1164 ( .A(n1515), .B(n1514), .CI(n1513), .CO(n1623), .S(n1468) );
  ADDFHX2 U1165 ( .A(n2607), .B(n2606), .CI(n2605), .CO(n2604), .S(n2964) );
  NOR2X1 U1166 ( .A(n4087), .B(n4086), .Y(n4509) );
  NOR2X1 U1167 ( .A(n3565), .B(n3564), .Y(n3570) );
  ADDFHX2 U1168 ( .A(n2227), .B(n2226), .CI(n2225), .CO(n2250), .S(n2246) );
  ADDFHX2 U1169 ( .A(n3189), .B(n3188), .CI(n3187), .CO(n3159), .S(n3190) );
  ADDFHX2 U1170 ( .A(n3230), .B(n3229), .CI(n3228), .CO(n3323), .S(n3322) );
  ADDFHX2 U1171 ( .A(n3048), .B(n3047), .CI(n3046), .CO(n3120), .S(n3158) );
  AND2XL U1172 ( .A(n3580), .B(n3579), .Y(n1117) );
  OAI21XL U1173 ( .A0(n2134), .A1(n2133), .B0(n2132), .Y(n1065) );
  ADDFHX2 U1174 ( .A(n1496), .B(n1495), .CI(n1494), .CO(n1571), .S(n1513) );
  NAND2BXL U1175 ( .AN(n3366), .B(n1110), .Y(n1109) );
  ADDFHX2 U1176 ( .A(n2819), .B(n2818), .CI(n2817), .CO(n2731), .S(n2820) );
  ADDFHX2 U1177 ( .A(n2867), .B(n2865), .CI(n2866), .CO(n2873), .S(n3337) );
  NAND2BXL U1178 ( .AN(n2549), .B(n1105), .Y(n1104) );
  ADDFHX2 U1179 ( .A(n3077), .B(n3076), .CI(n3075), .CO(n3153), .S(n3116) );
  ADDFHX2 U1180 ( .A(n2035), .B(n2034), .CI(n2033), .CO(n2142), .S(n2031) );
  ADDFHX2 U1181 ( .A(n2210), .B(n2209), .CI(n2208), .CO(n2247), .S(n2193) );
  ADDFHX2 U1182 ( .A(n2598), .B(n2597), .CI(n2596), .CO(n2605), .S(n2953) );
  ADDFX1 U1183 ( .A(n3555), .B(n3554), .CI(n3553), .CO(n3565), .S(n3549) );
  XOR3X2 U1184 ( .A(n2795), .B(n2793), .C(n2794), .Y(n2871) );
  NAND2XL U1185 ( .A(n1093), .B(n927), .Y(n1092) );
  ADDFHX2 U1186 ( .A(n1979), .B(n1978), .CI(n1977), .CO(n2033), .S(n1982) );
  ADDFX2 U1187 ( .A(n1613), .B(n1612), .CI(n1611), .CO(n1729), .S(n1615) );
  ADDFX1 U1188 ( .A(n2622), .B(n2621), .CI(n2620), .CO(n2611), .S(n2817) );
  ADDFHX2 U1189 ( .A(n1352), .B(n1351), .CI(n1350), .CO(n1496), .S(n1348) );
  ADDFHX2 U1190 ( .A(n2679), .B(n2678), .CI(n2677), .CO(n2683), .S(n2656) );
  ADDFHX2 U1191 ( .A(n2798), .B(n2797), .CI(n2796), .CO(n2816), .S(n2865) );
  ADDFHX2 U1192 ( .A(n2909), .B(n2908), .CI(n2907), .CO(n2922), .S(n3345) );
  NAND2BXL U1193 ( .AN(n3022), .B(n688), .Y(n687) );
  NAND2BXL U1194 ( .AN(n1936), .B(n1932), .Y(n1934) );
  OAI22X1 U1195 ( .A0(IN_VALID), .A1(n4648), .B0(n4664), .B1(n4647), .Y(A[9])
         );
  NAND2X1 U1196 ( .A(n985), .B(n984), .Y(n983) );
  ADDFHX2 U1197 ( .A(n3102), .B(n3101), .CI(n3100), .CO(n3142), .S(n3098) );
  NOR2X1 U1198 ( .A(n4091), .B(n4563), .Y(n4094) );
  NOR2X1 U1199 ( .A(n4091), .B(n4552), .Y(n3505) );
  NAND2BXL U1200 ( .AN(n3039), .B(n995), .Y(n994) );
  ADDFHX2 U1201 ( .A(n2577), .B(n2576), .CI(n2575), .CO(n2586), .S(n2609) );
  XOR2X1 U1202 ( .A(n2619), .B(n1051), .Y(n2628) );
  OAI22X1 U1203 ( .A0(IN_VALID), .A1(n4632), .B0(n4664), .B1(n4631), .Y(A[1])
         );
  OAI2BB1XL U1204 ( .A0N(n3446), .A1N(n3445), .B0(n2364), .Y(n3539) );
  OAI2BB1XL U1205 ( .A0N(n3450), .A1N(n3449), .B0(n3448), .Y(n3513) );
  ADDFHX2 U1206 ( .A(n2844), .B(n2843), .CI(n2842), .CO(n2853), .S(n2923) );
  OAI22X1 U1207 ( .A0(n4664), .A1(n3845), .B0(IN_VALID), .B1(n3844), .Y(A[6])
         );
  OAI2BB2X1 U1208 ( .B0(n1654), .B1(n1700), .A0N(n716), .A1N(n1173), .Y(n1722)
         );
  OAI2BB1X1 U1209 ( .A0N(n3112), .A1N(n3110), .B0(n1942), .Y(n1993) );
  OAI22X1 U1210 ( .A0(n1783), .A1(n1956), .B0(n1710), .B1(n1955), .Y(n1804) );
  INVX1 U1211 ( .A(n3011), .Y(n689) );
  OAI22X1 U1212 ( .A0(IN_VALID), .A1(n4637), .B0(n4664), .B1(n4636), .Y(A[8])
         );
  OAI2BB1X1 U1213 ( .A0N(n4111), .A1N(n4110), .B0(n4109), .Y(A[0]) );
  ADDHX1 U1214 ( .A(n2973), .B(n2972), .CO(n3038), .S(n2990) );
  NAND2XL U1215 ( .A(n895), .B(n894), .Y(n893) );
  INVXL U1216 ( .A(n3111), .Y(n987) );
  OAI22X1 U1217 ( .A0(n4664), .A1(n3833), .B0(IN_VALID), .B1(n3832), .Y(A[7])
         );
  OAI222X1 U1218 ( .A0(n1132), .A1(n3856), .B0(IN_VALID), .B1(n3850), .C0(
        n3849), .C1(n4664), .Y(A[3]) );
  OAI222X1 U1219 ( .A0(n3856), .A1(n4640), .B0(IN_VALID), .B1(n3855), .C0(
        n4664), .C1(n3854), .Y(A[4]) );
  OAI2BB1X1 U1220 ( .A0N(n3271), .A1N(n3269), .B0(n1480), .Y(n1562) );
  NAND2X1 U1221 ( .A(n728), .B(n734), .Y(n1886) );
  OAI211X1 U1222 ( .A0(IN_VALID), .A1(n3825), .B0(n3824), .C0(n3823), .Y(A[2])
         );
  OAI22X1 U1223 ( .A0(n4664), .A1(n3837), .B0(IN_VALID), .B1(n3836), .Y(A[5])
         );
  INVX1 U1224 ( .A(n1070), .Y(n2640) );
  NAND2BXL U1225 ( .AN(n2756), .B(n894), .Y(n892) );
  BUFX4 U1226 ( .A(n2849), .Y(n578) );
  NOR2X1 U1227 ( .A(n1124), .B(n4563), .Y(n2396) );
  INVX1 U1228 ( .A(n3487), .Y(n3489) );
  NOR2X1 U1229 ( .A(n1118), .B(n4563), .Y(n4495) );
  BUFX12 U1230 ( .A(n2022), .Y(n579) );
  OAI2BB1X1 U1231 ( .A0N(n4661), .A1N(in_out_cnt[10]), .B0(n4651), .Y(A[10])
         );
  BUFX12 U1232 ( .A(n3029), .Y(n580) );
  NOR2X1 U1233 ( .A(n4564), .B(n4552), .Y(n4557) );
  NOR2X1 U1234 ( .A(n4352), .B(n4552), .Y(n4346) );
  NOR2X1 U1235 ( .A(n4564), .B(n4563), .Y(n4571) );
  INVX1 U1236 ( .A(n4598), .Y(n4270) );
  XOR2XL U1237 ( .A(n4450), .B(n4449), .Y(n4496) );
  NOR2X1 U1238 ( .A(n4646), .B(n1131), .Y(n4634) );
  NOR2X1 U1239 ( .A(n4650), .B(n3829), .Y(n3822) );
  NOR2X1 U1240 ( .A(n4647), .B(n4660), .Y(n4667) );
  NAND2X1 U1241 ( .A(n3813), .B(rst_n), .Y(n3815) );
  NOR2X2 U1242 ( .A(n1281), .B(n643), .Y(n1186) );
  OAI211XL U1243 ( .A0(n4624), .A1(lay_cnt[1]), .B0(n672), .C0(n3852), .Y(
        n3826) );
  INVX1 U1244 ( .A(n2694), .Y(n2663) );
  OAI2BB1XL U1245 ( .A0N(n2755), .A1N(n2753), .B0(n657), .Y(n3444) );
  NAND2X1 U1246 ( .A(n3526), .B(n2102), .Y(n4563) );
  NAND2X1 U1247 ( .A(n3783), .B(rst_n), .Y(n3813) );
  INVXL U1248 ( .A(n3110), .Y(n581) );
  NOR2X1 U1249 ( .A(n3828), .B(is_row), .Y(n3831) );
  INVX1 U1250 ( .A(n3964), .Y(n3799) );
  OAI2BB1XL U1251 ( .A0N(n4078), .A1N(n4077), .B0(n4076), .Y(n4518) );
  OR2XL U1252 ( .A(n2127), .B(n2005), .Y(n637) );
  NOR2X1 U1253 ( .A(n4620), .B(is_row), .Y(n3841) );
  NAND2X1 U1254 ( .A(n3829), .B(n3858), .Y(n4502) );
  INVX1 U1255 ( .A(n3786), .Y(n4675) );
  NAND3X1 U1256 ( .A(n618), .B(n3812), .C(n3751), .Y(n3964) );
  INVX1 U1257 ( .A(n3776), .Y(n4102) );
  NOR2BX1 U1258 ( .AN(n3780), .B(n3637), .Y(n3786) );
  OR4X1 U1259 ( .A(n2073), .B(mode_val), .C(n604), .D(n3780), .Y(n2332) );
  INVX2 U1260 ( .A(n2940), .Y(n582) );
  NAND2X1 U1261 ( .A(n3776), .B(mode_val), .Y(n4234) );
  NOR2X1 U1262 ( .A(n2070), .B(n712), .Y(n3829) );
  NAND2X1 U1263 ( .A(n3798), .B(n2056), .Y(n2090) );
  INVX2 U1264 ( .A(n3112), .Y(n583) );
  BUFX8 U1265 ( .A(n1152), .Y(n3106) );
  BUFX8 U1266 ( .A(n1651), .Y(n2755) );
  OAI2BB1XL U1267 ( .A0N(butt_a_real[12]), .A1N(n4147), .B0(n4133), .Y(n529)
         );
  OAI2BB1XL U1268 ( .A0N(butt_a_imag[3]), .A1N(n4147), .B0(n4126), .Y(n543) );
  OAI2BB1XL U1269 ( .A0N(butt_a_real[11]), .A1N(n4147), .B0(n4134), .Y(n527)
         );
  XOR2X1 U1270 ( .A(n809), .B(n808), .Y(n807) );
  INVX2 U1271 ( .A(n2199), .Y(n584) );
  XOR3X2 U1272 ( .A(n2631), .B(n979), .C(n978), .Y(n3091) );
  NAND2X1 U1273 ( .A(n3784), .B(n2101), .Y(n3776) );
  XOR2X2 U1274 ( .A(n2464), .B(n2463), .Y(n2765) );
  INVX2 U1275 ( .A(n1173), .Y(n585) );
  OAI2BB1XL U1276 ( .A0N(butt_a_imag[2]), .A1N(n4147), .B0(n3996), .Y(n525) );
  XNOR3X2 U1277 ( .A(n1149), .B(n1158), .C(n1151), .Y(n1152) );
  OAI2BB1XL U1278 ( .A0N(butt_a_real[10]), .A1N(n4147), .B0(n4135), .Y(n523)
         );
  INVX2 U1279 ( .A(n1880), .Y(n586) );
  XOR2X2 U1280 ( .A(n1790), .B(n1789), .Y(n2362) );
  NOR2X1 U1281 ( .A(n3773), .B(n4640), .Y(n3810) );
  INVX2 U1282 ( .A(n1791), .Y(n587) );
  XNOR3X2 U1283 ( .A(n2433), .B(n2438), .C(n682), .Y(n2883) );
  XNOR3X2 U1284 ( .A(n1221), .B(n1226), .C(n1085), .Y(n1235) );
  NOR2X1 U1285 ( .A(n3837), .B(n4654), .Y(n4659) );
  XNOR2X2 U1286 ( .A(n1220), .B(n1228), .Y(n3173) );
  OAI2BB1XL U1287 ( .A0N(butt_b_real[4]), .A1N(n4186), .B0(n4162), .Y(n512) );
  NOR2X1 U1288 ( .A(n3816), .B(n712), .Y(n3846) );
  OAI2BB1XL U1289 ( .A0N(butt_b_real[12]), .A1N(n4186), .B0(n4154), .Y(n530)
         );
  NAND2X1 U1290 ( .A(n1222), .B(n1223), .Y(n1085) );
  OAI2BB1XL U1291 ( .A0N(butt_b_real[16]), .A1N(n4186), .B0(n4150), .Y(n538)
         );
  OAI2BB1XL U1292 ( .A0N(butt_b_real[6]), .A1N(n4186), .B0(n4160), .Y(n516) );
  INVX1 U1293 ( .A(n3028), .Y(n589) );
  OAI2BB1XL U1294 ( .A0N(butt_b_imag[8]), .A1N(n4186), .B0(n4176), .Y(n554) );
  NAND2X1 U1295 ( .A(n2750), .B(n2751), .Y(n978) );
  OAI2BB1XL U1296 ( .A0N(butt_b_real[17]), .A1N(n4186), .B0(n4149), .Y(n540)
         );
  XNOR2X2 U1297 ( .A(n2434), .B(n2435), .Y(n3084) );
  OAI2BB1XL U1298 ( .A0N(butt_b_real[10]), .A1N(n4186), .B0(n4156), .Y(n524)
         );
  OAI2BB1XL U1299 ( .A0N(butt_b_real[1]), .A1N(n4186), .B0(n4165), .Y(n506) );
  OAI2BB1XL U1300 ( .A0N(butt_b_imag[14]), .A1N(n4186), .B0(n4170), .Y(n492)
         );
  BUFX8 U1301 ( .A(n1340), .Y(n591) );
  NOR2X1 U1302 ( .A(n3847), .B(n4677), .Y(n3819) );
  OAI2BB1XL U1303 ( .A0N(butt_b_real[5]), .A1N(n4186), .B0(n4161), .Y(n514) );
  NOR2X1 U1304 ( .A(n4111), .B(n2081), .Y(n2082) );
  XOR2X2 U1305 ( .A(n2010), .B(n921), .Y(n920) );
  OAI2BB1XL U1306 ( .A0N(butt_b_real[14]), .A1N(n4186), .B0(n4152), .Y(n534)
         );
  XNOR3X2 U1307 ( .A(n668), .B(n1082), .C(n1083), .Y(n1079) );
  OAI2BB1XL U1308 ( .A0N(butt_b_real[7]), .A1N(n4186), .B0(n4159), .Y(n518) );
  OAI2BB1XL U1309 ( .A0N(butt_b_real[3]), .A1N(n4186), .B0(n4163), .Y(n510) );
  INVX2 U1310 ( .A(n3181), .Y(n593) );
  XNOR2X2 U1311 ( .A(n2469), .B(n2459), .Y(n2757) );
  OAI2BB1XL U1312 ( .A0N(butt_b_imag[13]), .A1N(n4186), .B0(n4171), .Y(n490)
         );
  NOR2X1 U1313 ( .A(n1211), .B(n2885), .Y(n1212) );
  OAI2BB1XL U1314 ( .A0N(butt_a_real[15]), .A1N(n4147), .B0(n4130), .Y(n535)
         );
  OAI2BB1XL U1315 ( .A0N(butt_a_imag[14]), .A1N(n4147), .B0(n4116), .Y(n491)
         );
  OAI2BB1XL U1316 ( .A0N(butt_a_imag[13]), .A1N(n4147), .B0(n4117), .Y(n489)
         );
  OAI2BB1XL U1317 ( .A0N(butt_a_imag[18]), .A1N(n4147), .B0(n4112), .Y(n499)
         );
  OAI2BB1XL U1318 ( .A0N(butt_a_imag[15]), .A1N(n4147), .B0(n4115), .Y(n493)
         );
  OAI2BB1XL U1319 ( .A0N(butt_a_imag[5]), .A1N(n4147), .B0(n4125), .Y(n547) );
  OAI2BB1XL U1320 ( .A0N(butt_a_real[1]), .A1N(n4147), .B0(n4144), .Y(n505) );
  OAI2BB1XL U1321 ( .A0N(butt_a_real[8]), .A1N(n4147), .B0(n4137), .Y(n519) );
  INVX2 U1322 ( .A(n3965), .Y(n605) );
  NOR2X1 U1323 ( .A(n2893), .B(n2885), .Y(n2894) );
  NOR2X1 U1324 ( .A(n2011), .B(n2010), .Y(n2012) );
  NOR2X1 U1325 ( .A(n2002), .B(n2411), .Y(n2003) );
  INVX1 U1326 ( .A(n922), .Y(n921) );
  OAI2BB1XL U1327 ( .A0N(butt_a_real[16]), .A1N(n4147), .B0(n4129), .Y(n537)
         );
  NAND2X1 U1328 ( .A(n1760), .B(n1759), .Y(n1765) );
  OAI2BB1XL U1329 ( .A0N(butt_a_imag[9]), .A1N(n4147), .B0(n4121), .Y(n555) );
  OAI2BB1XL U1330 ( .A0N(butt_a_imag[4]), .A1N(n4147), .B0(n3966), .Y(n545) );
  OAI2BB1XL U1331 ( .A0N(butt_a_real[17]), .A1N(n4147), .B0(n4128), .Y(n539)
         );
  NOR2X1 U1332 ( .A(n1635), .B(n2438), .Y(n1636) );
  NOR2X1 U1333 ( .A(n2411), .B(n2410), .Y(n2412) );
  NOR2X1 U1334 ( .A(n2080), .B(n2079), .Y(n2081) );
  NOR2X1 U1335 ( .A(n2439), .B(n2438), .Y(n2440) );
  NOR2X1 U1336 ( .A(n2001), .B(butt_b_real[17]), .Y(n1950) );
  NOR2X1 U1337 ( .A(Q[1]), .B(n2057), .Y(n3941) );
  NOR2X1 U1338 ( .A(n1892), .B(butt_a_imag[16]), .Y(n1016) );
  INVXL U1339 ( .A(n3867), .Y(n628) );
  NOR2X1 U1340 ( .A(n1331), .B(butt_b_real[7]), .Y(n1269) );
  NOR2X1 U1341 ( .A(n2409), .B(butt_a_real[17]), .Y(n2404) );
  NOR2X1 U1342 ( .A(n1251), .B(butt_a_imag[0]), .Y(n1250) );
  XOR2X2 U1343 ( .A(n1336), .B(butt_a_imag[8]), .Y(n1338) );
  NOR2X1 U1344 ( .A(n1196), .B(butt_b_real[5]), .Y(n1191) );
  NOR2X1 U1345 ( .A(n1180), .B(butt_b_real[3]), .Y(n1174) );
  NOR2X1 U1346 ( .A(n1210), .B(butt_b_real[1]), .Y(n1203) );
  NOR2X1 U1347 ( .A(n4104), .B(n4644), .Y(n3827) );
  NOR2X1 U1348 ( .A(n2437), .B(butt_a_real[11]), .Y(n2433) );
  NOR2X1 U1349 ( .A(n1767), .B(butt_a_imag[13]), .Y(n1646) );
  NOR2X1 U1350 ( .A(n1336), .B(butt_a_imag[8]), .Y(n1007) );
  NOR2X1 U1351 ( .A(n1751), .B(butt_b_real[13]), .Y(n909) );
  AND2X1 U1352 ( .A(lay_cnt[1]), .B(lay_cnt[0]), .Y(n3762) );
  INVX1 U1353 ( .A(in_out_cnt[3]), .Y(n3849) );
  INVX1 U1354 ( .A(lay_cnt[1]), .Y(n4104) );
  INVX1 U1355 ( .A(in_out_cnt[9]), .Y(n4647) );
  INVX1 U1356 ( .A(butt_b_imag[0]), .Y(n1251) );
  INVX1 U1357 ( .A(in_out_cnt[7]), .Y(n3833) );
  NOR2X1 U1358 ( .A(DP_OP_132J1_122_4436_n2999), .B(butt_a_real[0]), .Y(n2886)
         );
  BUFX2 U1359 ( .A(Q[16]), .Y(n3875) );
  INVX1 U1360 ( .A(in_out_cnt[5]), .Y(n3837) );
  NOR2X1 U1361 ( .A(Q[5]), .B(butt_a_imag[5]), .Y(n3668) );
  NOR2X1 U1362 ( .A(Q[31]), .B(butt_a_real[12]), .Y(n3497) );
  NOR2X1 U1363 ( .A(Q[3]), .B(butt_a_imag[3]), .Y(n4248) );
  OR2XL U1364 ( .A(Q[35]), .B(butt_a_real[16]), .Y(n3491) );
  NOR2X1 U1365 ( .A(Q[30]), .B(butt_a_real[11]), .Y(n4388) );
  NOR2X1 U1366 ( .A(Q[11]), .B(butt_a_imag[11]), .Y(n2389) );
  NOR2X1 U1367 ( .A(Q[29]), .B(butt_a_real[10]), .Y(n3729) );
  NOR2X1 U1368 ( .A(Q[9]), .B(butt_a_imag[9]), .Y(n3695) );
  NOR2X1 U1369 ( .A(Q[10]), .B(butt_a_imag[10]), .Y(n2088) );
  NOR2X1 U1370 ( .A(Q[28]), .B(butt_a_real[9]), .Y(n3731) );
  NOR2X1 U1371 ( .A(Q[27]), .B(butt_a_real[8]), .Y(n3736) );
  NOR2X1 U1372 ( .A(Q[22]), .B(butt_a_real[3]), .Y(n4277) );
  CLKBUFX1 U1373 ( .A(butt_b_real[11]), .Y(n681) );
  NOR2X1 U1374 ( .A(Q[21]), .B(butt_a_real[2]), .Y(n4275) );
  NOR2X1 U1375 ( .A(Q[20]), .B(butt_a_real[1]), .Y(n3910) );
  XOR2X2 U1376 ( .A(butt_b_imag[5]), .B(butt_a_imag[5]), .Y(n1228) );
  NOR2X1 U1377 ( .A(Q[13]), .B(butt_a_imag[13]), .Y(n4008) );
  XOR2X2 U1378 ( .A(butt_a_real[5]), .B(butt_b_real[5]), .Y(n2751) );
  OR2XL U1379 ( .A(Q[14]), .B(butt_a_imag[14]), .Y(n2075) );
  NOR2X1 U1380 ( .A(Q[15]), .B(butt_a_imag[15]), .Y(n2093) );
  OR2XL U1381 ( .A(Q[16]), .B(butt_a_imag[16]), .Y(n2382) );
  NOR2X1 U1382 ( .A(Q[12]), .B(butt_a_imag[12]), .Y(n4046) );
  XOR2X2 U1383 ( .A(butt_a_real[3]), .B(butt_b_real[3]), .Y(n2897) );
  MXI2X1 U1384 ( .A(n1353), .B(n1215), .S0(n1214), .Y(n1219) );
  INVXL U1385 ( .A(n2338), .Y(n595) );
  OAI22X1 U1386 ( .A0(n2861), .A1(n3087), .B0(n3085), .B1(n2927), .Y(n2920) );
  NAND4X1 U1387 ( .A(n4562), .B(n4561), .C(n4560), .D(n4559), .Y(D_imag[5]) );
  OAI22X2 U1388 ( .A0(n2901), .A1(n2940), .B0(n2938), .B1(n1997), .Y(n2935) );
  OAI21X1 U1389 ( .A0(n2872), .A1(n2871), .B0(n2873), .Y(n1066) );
  INVX2 U1390 ( .A(butt_b_real[13]), .Y(n2466) );
  INVX1 U1391 ( .A(n2902), .Y(n597) );
  NAND2X2 U1392 ( .A(n1025), .B(n3680), .Y(n1470) );
  OAI22X1 U1393 ( .A0(n2028), .A1(n2198), .B0(n2125), .B1(n2199), .Y(n2120) );
  OAI21X1 U1394 ( .A0(n1554), .A1(n1555), .B0(n1553), .Y(n671) );
  XOR2X1 U1395 ( .A(n3164), .B(n1045), .Y(n1044) );
  XNOR2X1 U1396 ( .A(n745), .B(n3237), .Y(n3257) );
  XOR2X1 U1397 ( .A(n1165), .B(butt_a_imag[2]), .Y(n1082) );
  OAI22X1 U1398 ( .A0(n2241), .A1(n2362), .B0(n2204), .B1(n2361), .Y(n2238) );
  XOR2X2 U1399 ( .A(n1036), .B(n575), .Y(n3005) );
  INVX4 U1400 ( .A(n1353), .Y(n832) );
  XNOR2X1 U1401 ( .A(n3451), .B(n3258), .Y(n3052) );
  OAI22X1 U1402 ( .A0(n3167), .A1(n3259), .B0(n3024), .B1(n3261), .Y(n3170) );
  NAND2BX2 U1403 ( .AN(n1282), .B(n1261), .Y(n1155) );
  INVX1 U1404 ( .A(n1261), .Y(n888) );
  OAI22X1 U1405 ( .A0(n3071), .A1(n3070), .B0(n3069), .B1(n3068), .Y(n3135) );
  OAI22X1 U1406 ( .A0(n1711), .A1(n2938), .B0(n1779), .B1(n2940), .Y(n1803) );
  ADDFHX4 U1407 ( .A(n1499), .B(n1498), .CI(n1497), .CO(n1549), .S(n1495) );
  XOR3X2 U1408 ( .A(n2904), .B(n2903), .C(n597), .Y(n3346) );
  NAND2X4 U1409 ( .A(n1608), .B(n1213), .Y(n1607) );
  OAI2BB1X2 U1410 ( .A0N(n1608), .A1N(n1607), .B0(n1606), .Y(n1642) );
  BUFX1 U1411 ( .A(n3649), .Y(n4033) );
  OAI2BB1X1 U1412 ( .A0N(n4594), .A1N(n4399), .B0(n3636), .Y(D_real[4]) );
  NAND2X2 U1413 ( .A(n3265), .B(n942), .Y(n941) );
  OAI21X1 U1414 ( .A0(n776), .A1(n3338), .B0(n3337), .Y(n775) );
  NAND2X4 U1415 ( .A(n2864), .B(n2863), .Y(n776) );
  NAND2BX2 U1416 ( .AN(n1353), .B(n1214), .Y(n948) );
  NAND2X1 U1417 ( .A(n1214), .B(n845), .Y(n1147) );
  NAND4X1 U1418 ( .A(n4577), .B(n4576), .C(n4575), .D(n4574), .Y(D_imag[6]) );
  ADDFHX4 U1419 ( .A(n3142), .B(n3141), .CI(n3140), .CO(n3383), .S(n3138) );
  INVX2 U1420 ( .A(n706), .Y(n4001) );
  OAI22X1 U1421 ( .A0(n2023), .A1(n2362), .B0(n1957), .B1(n2361), .Y(n2020) );
  XOR2X2 U1422 ( .A(n711), .B(n1120), .Y(n4491) );
  ADDHX1 U1423 ( .A(n2768), .B(n2767), .CO(n2800), .S(n2787) );
  NAND2X1 U1424 ( .A(n4532), .B(n4598), .Y(n3995) );
  NAND2X1 U1425 ( .A(n4532), .B(n4596), .Y(n4486) );
  OAI2BB1X2 U1426 ( .A0N(n4028), .A1N(n4000), .B0(n3999), .Y(n706) );
  NAND2X1 U1427 ( .A(n1934), .B(n1933), .Y(n1938) );
  OAI21X2 U1428 ( .A0(n1948), .A1(n1949), .B0(n1947), .Y(n749) );
  NOR2X1 U1429 ( .A(n2247), .B(n2248), .Y(n763) );
  NOR2BX2 U1430 ( .AN(n3270), .B(n3558), .Y(n1995) );
  OAI21X4 U1431 ( .A0(n1471), .A1(n3677), .B0(n1470), .Y(n3931) );
  AOI21X2 U1432 ( .A0(n1465), .A1(n4243), .B0(n1464), .Y(n3677) );
  NAND2XL U1433 ( .A(n673), .B(n1791), .Y(n1239) );
  NAND2X2 U1434 ( .A(n1285), .B(n1199), .Y(n1281) );
  OAI22X1 U1435 ( .A0(n1779), .A1(n2938), .B0(n1802), .B1(n2940), .Y(n1830) );
  OAI22X1 U1436 ( .A0(n1905), .A1(n2264), .B0(n2263), .B1(n1794), .Y(n1903) );
  XOR3X2 U1437 ( .A(n1904), .B(n865), .C(n1903), .Y(n1902) );
  INVX4 U1438 ( .A(n866), .Y(n865) );
  INVXL U1439 ( .A(n4433), .Y(n598) );
  INVX2 U1440 ( .A(n598), .Y(n599) );
  XNOR3X2 U1441 ( .A(n819), .B(n2109), .C(n2108), .Y(n2133) );
  NAND2X1 U1442 ( .A(n818), .B(n819), .Y(n817) );
  NAND2X1 U1443 ( .A(n1065), .B(n1064), .Y(n2183) );
  NAND2X2 U1444 ( .A(n3415), .B(n3416), .Y(n3714) );
  XNOR2X1 U1445 ( .A(n645), .B(n2711), .Y(n2578) );
  NAND2X2 U1446 ( .A(n3647), .B(n943), .Y(n1874) );
  ADDFHX1 U1447 ( .A(n1709), .B(n1708), .CI(n1707), .CO(n1842), .S(n1688) );
  MXI2X4 U1448 ( .A(n1284), .B(n1170), .S0(n1261), .Y(n2022) );
  NAND2X2 U1449 ( .A(n1866), .B(n1867), .Y(n3643) );
  OAI22X1 U1450 ( .A0(n645), .A1(n747), .B0(n2938), .B1(n1997), .Y(n1581) );
  AOI21XL U1451 ( .A0(n4432), .A1(n4614), .B0(n3708), .Y(n3709) );
  XNOR2X1 U1452 ( .A(n4036), .B(n3655), .Y(n4432) );
  INVX2 U1453 ( .A(butt_b_real[9]), .Y(n2424) );
  XOR2X2 U1454 ( .A(n2196), .B(n2186), .Y(n2187) );
  NAND2X1 U1455 ( .A(n601), .B(n889), .Y(n602) );
  NAND2X1 U1456 ( .A(n600), .B(n1113), .Y(n603) );
  NAND2X1 U1457 ( .A(n602), .B(n603), .Y(n4505) );
  INVXL U1458 ( .A(n1113), .Y(n601) );
  ADDFHX4 U1459 ( .A(n1923), .B(n1922), .CI(n1921), .CO(n1966), .S(n1927) );
  BUFX1 U1460 ( .A(n1258), .Y(n3818) );
  INVXL U1461 ( .A(n3779), .Y(n604) );
  NAND2X1 U1462 ( .A(n4505), .B(n4598), .Y(n4101) );
  INVXL U1463 ( .A(n4262), .Y(n606) );
  INVXL U1464 ( .A(n606), .Y(n607) );
  INVX1 U1465 ( .A(n1795), .Y(n608) );
  INVX2 U1466 ( .A(n608), .Y(n609) );
  OAI22X1 U1467 ( .A0(n1665), .A1(n3109), .B0(n1757), .B1(n3106), .Y(n1832) );
  AND2X1 U1468 ( .A(n3270), .B(n610), .Y(n2926) );
  INVXL U1469 ( .A(n2839), .Y(n610) );
  XNOR2X1 U1470 ( .A(n715), .B(n588), .Y(n3260) );
  OAI2BB2X2 U1471 ( .B0(n1956), .B1(n1505), .A0N(n612), .A1N(n611), .Y(n1492)
         );
  XOR2X1 U1472 ( .A(n3270), .B(n1954), .Y(n612) );
  XNOR2X1 U1473 ( .A(n3250), .B(n2711), .Y(n2579) );
  BUFX20 U1474 ( .A(n3006), .Y(n3250) );
  BUFX1 U1475 ( .A(n3370), .Y(n613) );
  OAI22X1 U1476 ( .A0(n2029), .A1(n3446), .B0(n1959), .B1(n3445), .Y(n2041) );
  XNOR2X1 U1477 ( .A(n3201), .B(n2567), .Y(n2029) );
  XNOR2X2 U1478 ( .A(n3270), .B(n2197), .Y(n1638) );
  ADDFHX4 U1479 ( .A(n1502), .B(n1501), .CI(n1500), .CO(n1548), .S(n1515) );
  NOR2X1 U1480 ( .A(n3320), .B(n3319), .Y(n3905) );
  ADDFHX1 U1481 ( .A(n3315), .B(n3314), .CI(n3313), .CO(n3321), .S(n3320) );
  XNOR2X1 U1482 ( .A(n3250), .B(n3258), .Y(n3262) );
  XNOR2X1 U1483 ( .A(n3014), .B(n2512), .Y(n2882) );
  XOR2X1 U1484 ( .A(n3014), .B(n3181), .Y(n859) );
  XOR2X1 U1485 ( .A(n3014), .B(n576), .Y(n986) );
  XNOR2X1 U1486 ( .A(n3014), .B(n657), .Y(n2117) );
  XNOR2X1 U1487 ( .A(n3014), .B(n2432), .Y(n2617) );
  XNOR2X2 U1488 ( .A(n579), .B(n1954), .Y(n1610) );
  OAI22X1 U1489 ( .A0(n3090), .A1(n3182), .B0(n3089), .B1(n3184), .Y(n3129) );
  OR2X1 U1490 ( .A(n3325), .B(n679), .Y(n614) );
  XNOR3X2 U1491 ( .A(n1781), .B(n874), .C(n1780), .Y(n1844) );
  AND2X2 U1492 ( .A(n3265), .B(n584), .Y(n1643) );
  ADDFHX1 U1493 ( .A(n2808), .B(n2807), .CI(n2806), .CO(n2952), .S(n2870) );
  XNOR3X2 U1494 ( .A(n3357), .B(n3355), .C(n2944), .Y(n3377) );
  OAI21X1 U1495 ( .A0(n1846), .A1(n1847), .B0(n1845), .Y(n1786) );
  OAI21X4 U1496 ( .A0(n2199), .A1(n609), .B0(n849), .Y(n848) );
  OAI2BB2X2 U1497 ( .B0(n2737), .B1(n2755), .A0N(n894), .A1N(n615), .Y(n2767)
         );
  INVX2 U1498 ( .A(n2753), .Y(n894) );
  OR2X2 U1499 ( .A(n1638), .B(n2198), .Y(n1639) );
  XNOR3X2 U1500 ( .A(n731), .B(n2603), .C(n2602), .Y(n616) );
  CLKINVX3 U1501 ( .A(n2604), .Y(n731) );
  ADDFHX4 U1502 ( .A(n1714), .B(n1712), .CI(n1713), .CO(n1813), .S(n1689) );
  ADDFHX1 U1503 ( .A(n2710), .B(n2709), .CI(n2708), .CO(n3437), .S(n2722) );
  NAND2X1 U1504 ( .A(n2910), .B(n3347), .Y(n2911) );
  XOR2X1 U1505 ( .A(n1074), .B(n2831), .Y(n2616) );
  OAI21X1 U1506 ( .A0(n2732), .A1(n1002), .B0(n2731), .Y(n868) );
  NAND2X1 U1507 ( .A(n4596), .B(n886), .Y(n4475) );
  XNOR2X1 U1508 ( .A(n3451), .B(n591), .Y(n1889) );
  XNOR2X1 U1509 ( .A(n3451), .B(n2432), .Y(n2473) );
  XOR3X4 U1510 ( .A(n3344), .B(n3343), .C(n3342), .Y(n3370) );
  NOR2BX2 U1511 ( .AN(n3270), .B(n4078), .Y(n2555) );
  NAND2X1 U1512 ( .A(n3998), .B(n2291), .Y(n2293) );
  AND2X2 U1513 ( .A(n3270), .B(n734), .Y(n1888) );
  INVXL U1514 ( .A(n2362), .Y(n734) );
  OAI2BB1X2 U1515 ( .A0N(n722), .A1N(n2048), .B0(n1056), .Y(n2140) );
  INVXL U1516 ( .A(n2048), .Y(n779) );
  XNOR2X1 U1517 ( .A(n3004), .B(n591), .Y(n1941) );
  XNOR2X1 U1518 ( .A(n769), .B(n3237), .Y(n1311) );
  BUFX1 U1519 ( .A(n4324), .Y(n721) );
  NAND2XL U1520 ( .A(n1640), .B(n1639), .Y(n1718) );
  XNOR2X1 U1521 ( .A(n3014), .B(n3237), .Y(n1237) );
  INVXL U1522 ( .A(n2361), .Y(n630) );
  OAI22X1 U1523 ( .A0(n2736), .A1(n2765), .B0(n2763), .B1(n977), .Y(n2768) );
  INVX1 U1524 ( .A(n1957), .Y(n728) );
  XNOR2X1 U1525 ( .A(n2783), .B(n1880), .Y(n1957) );
  NAND2X1 U1526 ( .A(n4460), .B(n3465), .Y(n3467) );
  OAI22X1 U1527 ( .A0(n2232), .A1(n2753), .B0(n2265), .B1(n2755), .Y(n2261) );
  XNOR2X1 U1528 ( .A(n2975), .B(n657), .Y(n2232) );
  NAND2X1 U1529 ( .A(n625), .B(n1095), .Y(n626) );
  XNOR2X1 U1530 ( .A(n3164), .B(n1791), .Y(n1602) );
  XNOR2X1 U1531 ( .A(n949), .B(n3173), .Y(n1543) );
  OAI22X1 U1532 ( .A0(n2672), .A1(n3450), .B0(n2539), .B1(n3449), .Y(n2679) );
  NAND2XL U1533 ( .A(n3336), .B(n3335), .Y(n617) );
  AOI21X1 U1534 ( .A0(n4595), .A1(n4598), .B0(n3710), .Y(n3711) );
  INVXL U1535 ( .A(n3778), .Y(n618) );
  AOI21X1 U1536 ( .A0(n3460), .A1(n3469), .B0(n3431), .Y(n3432) );
  BUFX12 U1537 ( .A(n1037), .Y(n1038) );
  NAND3X2 U1538 ( .A(n917), .B(n916), .C(n961), .Y(n1037) );
  XNOR2X1 U1539 ( .A(n1038), .B(n4076), .Y(n2487) );
  XNOR2X1 U1540 ( .A(n3164), .B(n1749), .Y(n2115) );
  OAI2BB1X4 U1541 ( .A0N(n762), .A1N(n2246), .B0(n761), .Y(n760) );
  INVX2 U1542 ( .A(n4578), .Y(n619) );
  NAND2BX1 U1543 ( .AN(n2917), .B(n767), .Y(n766) );
  OAI21X1 U1544 ( .A0(n2794), .A1(n2795), .B0(n2793), .Y(n2780) );
  ADDFHX4 U1545 ( .A(n2775), .B(n2774), .CI(n2773), .CO(n2795), .S(n2852) );
  OR2X4 U1546 ( .A(n913), .B(n3583), .Y(n804) );
  NAND2X1 U1547 ( .A(n840), .B(n1925), .Y(n839) );
  NAND2X4 U1548 ( .A(n2264), .B(n1754), .Y(n2263) );
  INVXL U1549 ( .A(n3239), .Y(n771) );
  NOR2BX1 U1550 ( .AN(n3239), .B(n3087), .Y(n3115) );
  XNOR2X1 U1551 ( .A(n3239), .B(n2432), .Y(n2847) );
  XNOR2X1 U1552 ( .A(n3239), .B(n591), .Y(n1356) );
  XNOR2X1 U1553 ( .A(n3239), .B(n2979), .Y(n1288) );
  XNOR2X1 U1554 ( .A(n3239), .B(n3084), .Y(n3086) );
  NAND2BX1 U1555 ( .AN(n3239), .B(n2757), .Y(n2736) );
  XNOR2X1 U1556 ( .A(n580), .B(n2979), .Y(n1544) );
  OAI2BB1X1 U1557 ( .A0N(n3106), .A1N(n3109), .B0(n1763), .Y(n1876) );
  NAND2BX2 U1558 ( .AN(n1857), .B(n1856), .Y(n1820) );
  BUFX2 U1559 ( .A(n3471), .Y(n3472) );
  XOR2X1 U1560 ( .A(n1038), .B(n657), .Y(n895) );
  XNOR2X2 U1561 ( .A(n2975), .B(n3237), .Y(n1525) );
  XNOR2X1 U1562 ( .A(n3265), .B(n1606), .Y(n1407) );
  XNOR2X1 U1563 ( .A(n3265), .B(n3253), .Y(n3255) );
  XNOR2X1 U1564 ( .A(n3265), .B(n1173), .Y(n1255) );
  OAI22X1 U1565 ( .A0(n3008), .A1(n3110), .B0(n1040), .B1(n3112), .Y(n3045) );
  XNOR2X1 U1566 ( .A(n3270), .B(n591), .Y(n3008) );
  ADDFHX4 U1567 ( .A(n1349), .B(n1348), .CI(n1347), .CO(n1514), .S(n1365) );
  AOI22X1 U1568 ( .A0(n620), .A1(n4598), .B0(n4589), .B1(n4594), .Y(n4577) );
  XNOR2X1 U1569 ( .A(n726), .B(n1880), .Y(n631) );
  INVXL U1570 ( .A(n2377), .Y(n2379) );
  INVX4 U1571 ( .A(n1240), .Y(n1284) );
  OAI2BB1X4 U1572 ( .A0N(n3998), .A1N(n2349), .B0(n4026), .Y(n778) );
  XOR2X2 U1573 ( .A(n4514), .B(n3458), .Y(n4097) );
  INVX1 U1574 ( .A(n4471), .Y(n3460) );
  NAND2X1 U1575 ( .A(n4522), .B(n622), .Y(n623) );
  NAND2X1 U1576 ( .A(n623), .B(n624), .Y(n4523) );
  CLKINVX2 U1577 ( .A(n4522), .Y(n621) );
  INVXL U1578 ( .A(n1119), .Y(n622) );
  XNOR2X1 U1579 ( .A(n3201), .B(n2432), .Y(n2829) );
  XNOR2X1 U1580 ( .A(n3201), .B(n2512), .Y(n3069) );
  XNOR2X1 U1581 ( .A(n3201), .B(n591), .Y(n1517) );
  XNOR2X1 U1582 ( .A(n3201), .B(n3173), .Y(n1295) );
  XNOR2X2 U1583 ( .A(n3201), .B(n2757), .Y(n2766) );
  OAI22XL U1584 ( .A0(n2792), .A1(n2883), .B0(n2846), .B1(n2829), .Y(n2796) );
  XOR2X2 U1585 ( .A(n579), .B(n1075), .Y(n1795) );
  NAND2X1 U1586 ( .A(n4228), .B(n4227), .Y(n4229) );
  OAI22X2 U1587 ( .A0(n1534), .A1(n2127), .B0(n2126), .B1(n2005), .Y(n1674) );
  NAND2X2 U1588 ( .A(n960), .B(n959), .Y(n885) );
  NAND2X4 U1589 ( .A(n726), .B(n772), .Y(n627) );
  BUFX8 U1590 ( .A(n3058), .Y(n1074) );
  ADDFHX4 U1591 ( .A(n2997), .B(n2996), .CI(n2995), .CO(n3002), .S(n3194) );
  BUFX8 U1592 ( .A(n3270), .Y(n3265) );
  MXI2X1 U1593 ( .A(n1280), .B(n1273), .S0(n764), .Y(n1187) );
  NAND2X1 U1594 ( .A(n3568), .B(n912), .Y(n834) );
  NAND2X1 U1595 ( .A(n912), .B(n911), .Y(n899) );
  NOR2X1 U1596 ( .A(n1995), .B(n1996), .Y(n819) );
  XNOR2X1 U1597 ( .A(n1995), .B(n1996), .Y(n2021) );
  XNOR3X2 U1598 ( .A(n731), .B(n2603), .C(n2602), .Y(n3422) );
  ADDFHX4 U1599 ( .A(n2583), .B(n2582), .CI(n2581), .CO(n2600), .S(n2653) );
  OAI22X2 U1600 ( .A0(n2838), .A1(n2839), .B0(n2837), .B1(n2836), .Y(n2904) );
  XOR3X2 U1601 ( .A(n3378), .B(n3379), .C(n3377), .Y(n880) );
  MXI2X2 U1602 ( .A(n845), .B(n1259), .S0(n844), .Y(n1164) );
  MXI2X2 U1603 ( .A(n1259), .B(n845), .S0(n897), .Y(n1260) );
  INVX8 U1604 ( .A(n1163), .Y(n845) );
  OAI22X1 U1605 ( .A0(n1774), .A1(n3110), .B0(n1889), .B1(n3112), .Y(n1875) );
  XOR2X1 U1606 ( .A(n971), .B(n1041), .Y(n1774) );
  OAI2BB2X2 U1607 ( .B0(n3868), .B1(n3866), .A0N(n628), .A1N(n570), .Y(
        FFT2D_OUT_R[0]) );
  NAND3X4 U1608 ( .A(n1208), .B(n1207), .C(n1206), .Y(n2733) );
  XNOR2X1 U1609 ( .A(n3164), .B(n657), .Y(n2444) );
  XNOR2X1 U1610 ( .A(n3054), .B(n657), .Y(n2490) );
  XNOR2X1 U1611 ( .A(n580), .B(n2512), .Y(n2931) );
  NAND3X4 U1612 ( .A(n1155), .B(n1216), .C(n1194), .Y(n3006) );
  OAI21X2 U1613 ( .A0(n3343), .A1(n3344), .B0(n3342), .Y(n2864) );
  OAI22X1 U1614 ( .A0(n1911), .A1(n2755), .B0(n1799), .B1(n2753), .Y(n1917) );
  BUFX8 U1615 ( .A(n1632), .Y(n2197) );
  INVX2 U1616 ( .A(n2197), .Y(n1075) );
  XNOR2X2 U1617 ( .A(n1888), .B(n1887), .Y(n1904) );
  NAND2X2 U1618 ( .A(n914), .B(n913), .Y(n912) );
  XOR2X1 U1619 ( .A(n627), .B(n1075), .Y(n1909) );
  OAI2BB1X2 U1620 ( .A0N(n4596), .A1N(n4578), .B0(n3709), .Y(n3710) );
  OAI2BB2X2 U1621 ( .B0(n3866), .B1(n3892), .A0N(n629), .A1N(n570), .Y(
        FFT2D_OUT_R[3]) );
  NAND2X4 U1622 ( .A(n3958), .B(n654), .Y(n4235) );
  OAI2BB1X2 U1623 ( .A0N(n630), .A1N(n631), .B0(n1886), .Y(n1935) );
  OAI211X1 U1624 ( .A0(n4321), .A1(n4541), .B0(n3634), .C0(n3633), .Y(n3635)
         );
  XNOR2X1 U1625 ( .A(n3004), .B(n2432), .Y(n2526) );
  XOR2X2 U1626 ( .A(n1250), .B(n1249), .Y(n1252) );
  INVX4 U1627 ( .A(n4459), .Y(n3967) );
  OAI2BB2X2 U1628 ( .B0(n3866), .B1(n3861), .A0N(n632), .A1N(n570), .Y(
        FFT2D_OUT_R[8]) );
  INVX4 U1629 ( .A(n1280), .Y(n1067) );
  XNOR2X2 U1630 ( .A(n1038), .B(n2830), .Y(n2784) );
  XNOR3X2 U1631 ( .A(n2822), .B(n1095), .C(n2820), .Y(n2950) );
  BUFX12 U1632 ( .A(n1148), .Y(n3201) );
  NAND4X1 U1633 ( .A(n4403), .B(n4402), .C(n4401), .D(n4400), .Y(D_real[9]) );
  NAND4X1 U1634 ( .A(n4414), .B(n4412), .C(n4413), .D(n4411), .Y(D_real[10])
         );
  ADDFHX4 U1635 ( .A(n2856), .B(n2855), .CI(n2854), .CO(n2875), .S(n3343) );
  NAND2X1 U1636 ( .A(n4485), .B(n4596), .Y(n4413) );
  NAND2X4 U1637 ( .A(n770), .B(n1194), .Y(n750) );
  OAI2BB2X2 U1638 ( .B0(n3866), .B1(n3878), .A0N(n633), .A1N(n570), .Y(
        FFT2D_OUT_R[9]) );
  NAND2X1 U1639 ( .A(n3998), .B(n2322), .Y(n2324) );
  INVX4 U1640 ( .A(n4024), .Y(n3998) );
  OAI22X1 U1641 ( .A0(n2114), .A1(n3558), .B0(n2004), .B1(n3557), .Y(n2108) );
  XNOR2X1 U1642 ( .A(n3270), .B(n3556), .Y(n2004) );
  NAND2X1 U1643 ( .A(n2000), .B(n1999), .Y(n3542) );
  OAI21X2 U1644 ( .A0(n4514), .A1(n3508), .B0(n4069), .Y(n791) );
  OAI21X2 U1645 ( .A0(n3471), .A1(n935), .B0(n931), .Y(n930) );
  BUFX8 U1646 ( .A(n1503), .Y(n3451) );
  INVX4 U1647 ( .A(n2349), .Y(n4027) );
  NAND2X2 U1648 ( .A(n2349), .B(n2348), .Y(n913) );
  ADDFHX1 U1649 ( .A(n1361), .B(n1360), .CI(n1359), .CO(n1497), .S(n1364) );
  XNOR2X1 U1650 ( .A(n1036), .B(n2979), .Y(n2826) );
  OAI22X1 U1651 ( .A0(n2905), .A1(n3109), .B0(n3106), .B1(n2826), .Y(n2879) );
  OAI22X1 U1652 ( .A0(n1542), .A1(n2938), .B0(n1609), .B1(n2940), .Y(n1590) );
  XNOR2X1 U1653 ( .A(n3250), .B(n2900), .Y(n1609) );
  OAI211X1 U1654 ( .A0(n4551), .A1(n4541), .B0(n3684), .C0(n3683), .Y(n3685)
         );
  INVX2 U1655 ( .A(n1185), .Y(n1194) );
  XOR3X2 U1656 ( .A(n3039), .B(n996), .C(n3038), .Y(n3033) );
  OAI2BB1X4 U1657 ( .A0N(n4460), .A1N(n4469), .B0(n3472), .Y(n854) );
  NAND2X2 U1658 ( .A(n945), .B(n941), .Y(n944) );
  INVX2 U1659 ( .A(n3471), .Y(n4467) );
  AOI21X1 U1660 ( .A0(n4596), .A1(n4491), .B0(n3507), .Y(n3525) );
  NAND2X1 U1661 ( .A(n746), .B(n3506), .Y(n3507) );
  INVX2 U1662 ( .A(cs[0]), .Y(n3750) );
  XNOR2X1 U1663 ( .A(n3451), .B(n2830), .Y(n2161) );
  NAND4X1 U1664 ( .A(n4478), .B(n4477), .C(n4476), .D(n4475), .Y(D_real[13])
         );
  OAI21X1 U1665 ( .A0(n2869), .A1(n2870), .B0(n2868), .Y(n2805) );
  NAND2BX2 U1666 ( .AN(n4292), .B(n4272), .Y(n680) );
  NAND3X1 U1667 ( .A(n1276), .B(n1142), .C(n947), .Y(n946) );
  NAND2X1 U1668 ( .A(n1276), .B(n1353), .Y(n1277) );
  NAND2X1 U1669 ( .A(cs[2]), .B(cs[0]), .Y(n1011) );
  MXI2X1 U1670 ( .A(lay_cnt[3]), .B(lay_cnt[2]), .S0(cs[0]), .Y(n1134) );
  OAI21X2 U1671 ( .A0(n4379), .A1(n3971), .B0(n3970), .Y(n3973) );
  OAI22X1 U1672 ( .A0(n2556), .A1(n2753), .B0(n2444), .B1(n2755), .Y(n2559) );
  NAND2X2 U1673 ( .A(n1198), .B(n1282), .Y(n1208) );
  NAND2X4 U1674 ( .A(n1231), .B(n1162), .Y(n1282) );
  INVX4 U1675 ( .A(n1184), .Y(n1136) );
  AOI21X4 U1676 ( .A0(n933), .A1(n4469), .B0(n930), .Y(n4514) );
  NAND2X1 U1677 ( .A(n4504), .B(n4596), .Y(n4536) );
  XNOR2X1 U1678 ( .A(n3250), .B(n2674), .Y(n2458) );
  OAI21X1 U1679 ( .A0(n4514), .A1(n4506), .B0(n4510), .Y(n889) );
  NOR2X1 U1680 ( .A(n1231), .B(n1167), .Y(n1185) );
  ADDFHX1 U1681 ( .A(n2693), .B(n2692), .CI(n2694), .CO(n2710), .S(n2689) );
  XOR2XL U1682 ( .A(n2437), .B(n2436), .Y(n2439) );
  XOR2XL U1683 ( .A(n1634), .B(n1633), .Y(n1635) );
  NOR2X1 U1684 ( .A(n1531), .B(n2425), .Y(n1532) );
  NAND2X1 U1685 ( .A(n1270), .B(n2639), .Y(n869) );
  XNOR2X1 U1686 ( .A(n2746), .B(n1174), .Y(n1178) );
  NAND2X1 U1687 ( .A(n1192), .B(n2751), .Y(n952) );
  NOR2X1 U1688 ( .A(n1883), .B(n733), .Y(n1884) );
  OAI21XL U1689 ( .A0(n4012), .A1(n4008), .B0(n4009), .Y(n2077) );
  NAND2X1 U1690 ( .A(n2434), .B(n2435), .Y(n682) );
  OR2XL U1691 ( .A(n1166), .B(n2057), .Y(n668) );
  XOR2XL U1692 ( .A(n871), .B(n2511), .Y(n870) );
  NOR2X1 U1693 ( .A(n1332), .B(n2506), .Y(n871) );
  INVXL U1694 ( .A(n1338), .Y(n810) );
  NOR2X1 U1695 ( .A(n1181), .B(n2746), .Y(n1182) );
  XOR2XL U1696 ( .A(n1180), .B(n1179), .Y(n1181) );
  XOR2X1 U1697 ( .A(n955), .B(n954), .Y(n953) );
  INVXL U1698 ( .A(n2639), .Y(n954) );
  NAND2X1 U1699 ( .A(n2469), .B(n2459), .Y(n2449) );
  OAI22XL U1700 ( .A0(n2738), .A1(n2836), .B0(n2616), .B1(n2839), .Y(n2802) );
  NAND2X1 U1701 ( .A(n890), .B(n892), .Y(n2803) );
  BUFX3 U1702 ( .A(n3360), .Y(n727) );
  INVX2 U1703 ( .A(n1069), .Y(n1068) );
  NOR2X1 U1704 ( .A(n2636), .B(n2632), .Y(n2637) );
  XOR2X1 U1705 ( .A(n1225), .B(n1224), .Y(n1227) );
  OAI22XL U1706 ( .A0(n2305), .A1(n4078), .B0(n2270), .B1(n4077), .Y(n2302) );
  OAI22XL U1707 ( .A0(n2268), .A1(n2361), .B0(n2301), .B1(n2362), .Y(n2304) );
  NOR2X1 U1708 ( .A(n2178), .B(n3557), .Y(n828) );
  NAND2BXL U1709 ( .AN(n819), .B(n2109), .Y(n816) );
  OAI22XL U1710 ( .A0(n1973), .A1(n2755), .B0(n2753), .B1(n1911), .Y(n1962) );
  OAI22XL U1711 ( .A0(n1909), .A1(n2198), .B0(n1972), .B1(n2199), .Y(n1964) );
  OAI22XL U1712 ( .A0(n3543), .A1(n3557), .B0(n3558), .B1(n3542), .Y(n3561) );
  NAND2XL U1713 ( .A(n3548), .B(n3585), .Y(n3567) );
  AOI21XL U1714 ( .A0(n2083), .A1(n2067), .B0(n2066), .Y(n4012) );
  NOR2X1 U1715 ( .A(n4044), .B(n4046), .Y(n2067) );
  INVXL U1716 ( .A(n2083), .Y(n4045) );
  XNOR2X1 U1717 ( .A(n3234), .B(n2711), .Y(n2472) );
  INVX2 U1718 ( .A(n2900), .Y(n1997) );
  XNOR2X1 U1719 ( .A(n3054), .B(n591), .Y(n2827) );
  XOR2X1 U1720 ( .A(n579), .B(n591), .Y(n990) );
  XNOR2XL U1721 ( .A(n579), .B(n2979), .Y(n3059) );
  XNOR2X1 U1722 ( .A(n769), .B(n3028), .Y(n3030) );
  XNOR2XL U1723 ( .A(n949), .B(n657), .Y(n2177) );
  AND2X1 U1724 ( .A(n1699), .B(n2462), .Y(n910) );
  XOR2X1 U1725 ( .A(n2467), .B(n909), .Y(n908) );
  XOR2XL U1726 ( .A(n1753), .B(n2469), .Y(n1754) );
  NOR2X1 U1727 ( .A(n1752), .B(n2467), .Y(n1753) );
  XOR2XL U1728 ( .A(n1751), .B(n1750), .Y(n1752) );
  ADDHXL U1729 ( .A(n1293), .B(n1292), .CO(n1266), .S(n1309) );
  NOR2BX1 U1730 ( .AN(n3270), .B(n1793), .Y(n1293) );
  NOR2BX1 U1731 ( .AN(n645), .B(n3106), .Y(n1292) );
  NAND2XL U1732 ( .A(butt_b_real[18]), .B(n4673), .Y(n2402) );
  OAI21XL U1733 ( .A0(butt_b_real[18]), .A1(n4673), .B0(butt_a_real[17]), .Y(
        n2403) );
  NAND2XL U1734 ( .A(butt_b_imag[18]), .B(n3530), .Y(n2007) );
  OAI21XL U1735 ( .A0(butt_b_imag[18]), .A1(n3530), .B0(butt_a_imag[17]), .Y(
        n2008) );
  OAI2BB1XL U1736 ( .A0N(n3446), .A1N(n3445), .B0(n2567), .Y(n4085) );
  XNOR2XL U1737 ( .A(n580), .B(n2711), .Y(n2491) );
  OAI22XL U1738 ( .A0(n3446), .A1(n2498), .B0(n3445), .B1(n1014), .Y(n2560) );
  OAI22XL U1739 ( .A0(n2595), .A1(n2763), .B0(n2565), .B1(n2765), .Y(n2623) );
  OAI22XL U1740 ( .A0(n2766), .A1(n2765), .B0(n2764), .B1(n2763), .Y(n2801) );
  OAI22XL U1741 ( .A0(n2792), .A1(n2846), .B0(n2735), .B1(n2883), .Y(n2760) );
  OAI22X1 U1742 ( .A0(n2734), .A1(n2940), .B0(n2790), .B1(n2938), .Y(n2761) );
  NAND2X1 U1743 ( .A(n1098), .B(n1096), .Y(n2762) );
  INVX2 U1744 ( .A(n3372), .Y(n937) );
  OAI2BB1X1 U1745 ( .A0N(n3184), .A1N(n3182), .B0(n2752), .Y(n2843) );
  NAND2X1 U1746 ( .A(n847), .B(n846), .Y(n1922) );
  OAI22XL U1747 ( .A0(n1973), .A1(n2753), .B0(n2026), .B1(n2755), .Y(n2036) );
  OAI22XL U1748 ( .A0(n1899), .A1(n2938), .B0(n1943), .B1(n2940), .Y(n1944) );
  NAND2XL U1749 ( .A(n1936), .B(n1935), .Y(n1937) );
  OAI22XL U1750 ( .A0(n2128), .A1(n2362), .B0(n2023), .B1(n2361), .Y(n2131) );
  OAI22XL U1751 ( .A0(n2026), .A1(n2753), .B0(n2117), .B1(n2755), .Y(n2129) );
  OAI22XL U1752 ( .A0(n2014), .A1(n2839), .B0(n1961), .B1(n2836), .Y(n2039) );
  AND2X2 U1753 ( .A(n1960), .B(n919), .Y(n2040) );
  OAI22XL U1754 ( .A0(n1253), .A1(n1701), .B0(n1700), .B1(n585), .Y(n1373) );
  XOR2XL U1755 ( .A(n1212), .B(n2897), .Y(n1213) );
  NOR2BXL U1756 ( .AN(n3270), .B(n1608), .Y(n1405) );
  OAI22XL U1757 ( .A0(n1543), .A1(n3179), .B0(n1472), .B1(n3177), .Y(n1566) );
  OAI22X1 U1758 ( .A0(n1326), .A1(n3177), .B0(n1472), .B1(n3179), .Y(n1486) );
  NOR2X1 U1759 ( .A(n3661), .B(n3668), .Y(n3658) );
  NAND2X2 U1760 ( .A(n749), .B(n748), .Y(n2048) );
  NOR2X1 U1761 ( .A(Q[4]), .B(butt_a_imag[4]), .Y(n3661) );
  AOI21XL U1762 ( .A0(n2059), .A1(n3946), .B0(n2058), .Y(n3656) );
  NOR2X1 U1763 ( .A(n4246), .B(n4248), .Y(n2059) );
  NAND2X1 U1764 ( .A(n675), .B(n674), .Y(n1812) );
  XOR2XL U1765 ( .A(n1017), .B(n2413), .Y(n4079) );
  NAND2X1 U1766 ( .A(n2667), .B(n2668), .Y(n906) );
  OAI21X1 U1767 ( .A0(n2667), .A1(n2668), .B0(n2666), .Y(n907) );
  XOR3X2 U1768 ( .A(n2531), .B(n983), .C(n2532), .Y(n2534) );
  NAND2XL U1769 ( .A(n1744), .B(n1746), .Y(n723) );
  OAI21XL U1770 ( .A0(n3618), .A1(n3614), .B0(n3619), .Y(n3607) );
  NOR2X1 U1771 ( .A(n3611), .B(n3618), .Y(n3608) );
  OAI21XL U1772 ( .A0(n3357), .A1(n3356), .B0(n3355), .Y(n2942) );
  NAND2XL U1773 ( .A(n2772), .B(n2771), .Y(n1008) );
  NAND2BXL U1774 ( .AN(n2772), .B(n684), .Y(n683) );
  XOR3X2 U1775 ( .A(n2626), .B(n2627), .C(n2628), .Y(n2818) );
  NOR2X1 U1776 ( .A(n3288), .B(n3287), .Y(n3286) );
  INVXL U1777 ( .A(n3563), .Y(n3540) );
  OAI22XL U1778 ( .A0(n2365), .A1(n4077), .B0(n3541), .B1(n4078), .Y(n3538) );
  NAND2XL U1779 ( .A(n2247), .B(n2248), .Y(n761) );
  NAND2BX1 U1780 ( .AN(n2193), .B(n813), .Y(n812) );
  INVXL U1781 ( .A(n2194), .Y(n813) );
  NAND2XL U1782 ( .A(n2194), .B(n2193), .Y(n2195) );
  INVXL U1783 ( .A(n3656), .Y(n3667) );
  NAND2XL U1784 ( .A(Q[25]), .B(butt_a_real[6]), .Y(n4334) );
  AOI21XL U1785 ( .A0(n3617), .A1(n3608), .B0(n3607), .Y(n4336) );
  INVXL U1786 ( .A(n3494), .Y(n3740) );
  INVXL U1787 ( .A(n3606), .Y(n3617) );
  NAND2XL U1788 ( .A(n3160), .B(n3159), .Y(n707) );
  INVXL U1789 ( .A(n3160), .Y(n709) );
  NAND2X1 U1790 ( .A(n1939), .B(n1940), .Y(n923) );
  INVXL U1791 ( .A(n2098), .Y(n3526) );
  XOR3X2 U1792 ( .A(n2250), .B(n760), .C(n2249), .Y(n2283) );
  OAI21XL U1793 ( .A0(n4045), .A1(n2087), .B0(n2086), .Y(n2388) );
  AOI22XL U1794 ( .A0(n4608), .A1(FFT2D_IN_R[9]), .B0(n4607), .B1(n4606), .Y(
        n4609) );
  XOR2XL U1795 ( .A(n4045), .B(n3703), .Y(n4580) );
  OAI21XL U1796 ( .A0(n4464), .A1(n3463), .B0(n3462), .Y(n3464) );
  OAI2BB1XL U1797 ( .A0N(n3829), .A1N(n3526), .B0(n4563), .Y(n4530) );
  INVXL U1798 ( .A(n3567), .Y(n911) );
  AOI21X1 U1799 ( .A0(n3552), .A1(n3585), .B0(n3551), .Y(n3571) );
  XNOR2XL U1800 ( .A(n2077), .B(n2076), .Y(n4208) );
  XOR2XL U1801 ( .A(n4012), .B(n4011), .Y(n4207) );
  XNOR2XL U1802 ( .A(n4050), .B(n4049), .Y(n4221) );
  BUFX1 U1803 ( .A(n3752), .Y(n3806) );
  AOI21XL U1804 ( .A0(n4441), .A1(n4614), .B0(n4440), .Y(n4442) );
  NAND4XL U1805 ( .A(n4439), .B(n4438), .C(n4437), .D(n4436), .Y(n4440) );
  AOI21XL U1806 ( .A0(n4410), .A1(n4614), .B0(n4409), .Y(n4411) );
  NAND4XL U1807 ( .A(n4408), .B(n4407), .C(n4406), .D(n4405), .Y(n4409) );
  AOI21XL U1808 ( .A0(n4399), .A1(n4614), .B0(n4398), .Y(n4400) );
  NAND4XL U1809 ( .A(n4397), .B(n4396), .C(n4395), .D(n4394), .Y(n4398) );
  XOR2X1 U1810 ( .A(n1036), .B(n591), .Y(n1097) );
  INVX2 U1811 ( .A(n3173), .Y(n1045) );
  NAND2X1 U1812 ( .A(n1792), .B(n1793), .Y(n951) );
  XNOR2XL U1813 ( .A(n3004), .B(n2979), .Y(n1762) );
  XNOR2X1 U1814 ( .A(n1038), .B(n2197), .Y(n1778) );
  XNOR2XL U1815 ( .A(n645), .B(n2900), .Y(n1542) );
  XOR2X2 U1816 ( .A(n2975), .B(n1045), .Y(n1087) );
  XOR2X1 U1817 ( .A(n971), .B(n976), .Y(n2442) );
  XOR2X1 U1818 ( .A(n627), .B(n592), .Y(n2556) );
  INVX2 U1819 ( .A(n2555), .Y(n699) );
  NAND2X1 U1820 ( .A(n806), .B(n591), .Y(n2554) );
  NAND2XL U1821 ( .A(n3110), .B(n3112), .Y(n806) );
  XNOR2X1 U1822 ( .A(n1038), .B(n2567), .Y(n1014) );
  NAND2XL U1823 ( .A(n1097), .B(n581), .Y(n701) );
  NAND2XL U1824 ( .A(n591), .B(n583), .Y(n700) );
  INVXL U1825 ( .A(n3084), .Y(n974) );
  XNOR2X1 U1826 ( .A(n3004), .B(n2512), .Y(n2572) );
  XNOR2XL U1827 ( .A(n579), .B(n657), .Y(n2618) );
  OAI2BB1X1 U1828 ( .A0N(n3106), .A1N(n3109), .B0(n2979), .Y(n2614) );
  NAND2BX1 U1829 ( .AN(n3270), .B(n657), .Y(n2737) );
  XNOR2X1 U1830 ( .A(n949), .B(n2512), .Y(n2834) );
  XNOR2X1 U1831 ( .A(n3250), .B(n2432), .Y(n2848) );
  XNOR2X1 U1832 ( .A(n3270), .B(n2979), .Y(n2982) );
  XNOR2X1 U1833 ( .A(n1038), .B(n2979), .Y(n2967) );
  NAND2BXL U1834 ( .AN(n3270), .B(n591), .Y(n2969) );
  NAND2BX1 U1835 ( .AN(n3239), .B(n2512), .Y(n2970) );
  XNOR2XL U1836 ( .A(n1038), .B(n1749), .Y(n1905) );
  OAI22X1 U1837 ( .A0(n1777), .A1(n2755), .B0(n2753), .B1(n592), .Y(n1800) );
  NAND2BXL U1838 ( .AN(n645), .B(n657), .Y(n1777) );
  OAI22X1 U1839 ( .A0(n1671), .A1(n2839), .B0(n2836), .B1(n2831), .Y(n1704) );
  XNOR2XL U1840 ( .A(n3164), .B(n1880), .Y(n2204) );
  OAI22XL U1841 ( .A0(n2161), .A1(n2836), .B0(n2200), .B1(n2839), .Y(n2218) );
  OAI22XL U1842 ( .A0(n2164), .A1(n2198), .B0(n2199), .B1(n1075), .Y(n2216) );
  XNOR2XL U1843 ( .A(n1038), .B(n1880), .Y(n2023) );
  XOR2XL U1844 ( .A(n627), .B(n697), .Y(n2027) );
  OAI22X2 U1845 ( .A0(n1907), .A1(n3446), .B0(n901), .B1(n3445), .Y(n919) );
  NAND2BX1 U1846 ( .AN(n3239), .B(n2567), .Y(n1907) );
  XOR2XL U1847 ( .A(n1074), .B(n1539), .Y(n1245) );
  OAI22X1 U1848 ( .A0(n1241), .A1(n3106), .B0(n3109), .B1(n669), .Y(n1267) );
  XNOR2XL U1849 ( .A(n3166), .B(n591), .Y(n1593) );
  XNOR2X1 U1850 ( .A(n1037), .B(n1954), .Y(n1560) );
  XNOR2X1 U1851 ( .A(n3054), .B(n1173), .Y(n1516) );
  OAI2BB1X2 U1852 ( .A0N(n873), .A1N(n1780), .B0(n872), .Y(n1847) );
  INVXL U1853 ( .A(n1781), .Y(n875) );
  NOR2BXL U1854 ( .AN(n645), .B(n2755), .Y(n1834) );
  OAI2BB1X1 U1855 ( .A0N(n3179), .A1N(n3177), .B0(n1653), .Y(n1833) );
  INVXL U1856 ( .A(n853), .Y(n852) );
  OAI22XL U1857 ( .A0(n1711), .A1(n2940), .B0(n1678), .B1(n2938), .Y(n1708) );
  OAI22X2 U1858 ( .A0(n1591), .A1(n3109), .B0(n1666), .B1(n3106), .Y(n853) );
  OAI22XL U1859 ( .A0(n1678), .A1(n2940), .B0(n1609), .B1(n2938), .Y(n1681) );
  OAI2BB1X1 U1860 ( .A0N(n2765), .A1N(n2763), .B0(n2696), .Y(n2720) );
  OAI22XL U1861 ( .A0(n2713), .A1(n3445), .B0(n3446), .B1(n901), .Y(n3442) );
  OAI22XL U1862 ( .A0(n2712), .A1(n3449), .B0(n3447), .B1(n3450), .Y(n3443) );
  XNOR2XL U1863 ( .A(n2976), .B(n657), .Y(n2529) );
  XOR2X1 U1864 ( .A(n1074), .B(n901), .Y(n2489) );
  XNOR2X1 U1865 ( .A(n2675), .B(n2711), .Y(n2539) );
  OAI22XL U1866 ( .A0(n2472), .A1(n3449), .B0(n2491), .B1(n3450), .Y(n2483) );
  OAI22XL U1867 ( .A0(n2756), .A1(n2755), .B0(n2754), .B1(n2753), .Y(n2773) );
  OAI22X1 U1868 ( .A0(n2827), .A1(n3110), .B0(n2789), .B1(n3112), .Y(n2798) );
  OAI22X1 U1869 ( .A0(n2784), .A1(n2839), .B0(n2836), .B1(n2838), .Y(n2858) );
  XNOR2X1 U1870 ( .A(n3270), .B(n2830), .Y(n2837) );
  NAND2X1 U1871 ( .A(n881), .B(n3253), .Y(n2925) );
  NAND2XL U1872 ( .A(n3256), .B(n3254), .Y(n881) );
  XNOR2XL U1873 ( .A(n3250), .B(n3084), .Y(n3088) );
  XNOR2XL U1874 ( .A(n769), .B(n2512), .Y(n3071) );
  OAI22XL U1875 ( .A0(n2928), .A1(n3110), .B0(n2862), .B1(n3112), .Y(n2919) );
  OAI2BB1X1 U1876 ( .A0N(n987), .A1N(n581), .B0(n988), .Y(n3150) );
  OAI22XL U1877 ( .A0(n3059), .A1(n3109), .B0(n3108), .B1(n3106), .Y(n3100) );
  OAI22X1 U1878 ( .A0(n1084), .A1(n3256), .B0(n3254), .B1(n3055), .Y(n3102) );
  XNOR2XL U1879 ( .A(n949), .B(n594), .Y(n1263) );
  OAI22XL U1880 ( .A0(n3174), .A1(n3179), .B0(n3177), .B1(n1045), .Y(n3214) );
  XOR2XL U1881 ( .A(n2892), .B(n2891), .Y(n2893) );
  OAI22X1 U1882 ( .A0(n3090), .A1(n3184), .B0(n856), .B1(n3182), .Y(n3105) );
  XNOR2XL U1883 ( .A(n580), .B(n4076), .Y(n2240) );
  OAI22XL U1884 ( .A0(n2301), .A1(n2361), .B0(n2362), .B1(n586), .Y(n2357) );
  OAI22XL U1885 ( .A0(n2300), .A1(n3445), .B0(n2363), .B1(n3446), .Y(n2358) );
  INVXL U1886 ( .A(n2359), .Y(n2309) );
  OAI22XL U1887 ( .A0(n2267), .A1(n3445), .B0(n2300), .B1(n3446), .Y(n2307) );
  OAI22XL U1888 ( .A0(n2233), .A1(n2263), .B0(n2264), .B1(n697), .Y(n2260) );
  OAI22X1 U1889 ( .A0(n2177), .A1(n2755), .B0(n2753), .B1(n2117), .Y(n2175) );
  OAI22XL U1890 ( .A0(n2179), .A1(n4078), .B0(n2116), .B1(n4077), .Y(n2176) );
  OAI22X1 U1891 ( .A0(n2177), .A1(n2753), .B0(n2202), .B1(n2755), .Y(n2207) );
  OAI22XL U1892 ( .A0(n2202), .A1(n2753), .B0(n2232), .B1(n2755), .Y(n2229) );
  OAI22XL U1893 ( .A0(n1394), .A1(n3273), .B0(n1257), .B1(n3275), .Y(n1378) );
  NOR2BX1 U1894 ( .AN(n3270), .B(n1701), .Y(n1375) );
  XOR2X1 U1895 ( .A(n1223), .B(n1081), .Y(n1080) );
  INVX2 U1896 ( .A(n1079), .Y(n882) );
  NOR2X1 U1897 ( .A(n1078), .B(n1082), .Y(n1081) );
  OAI22XL U1898 ( .A0(n1264), .A1(n3177), .B0(n1326), .B1(n3179), .Y(n1319) );
  OAI22X1 U1899 ( .A0(n1324), .A1(n1793), .B0(n1792), .B1(n1287), .Y(n1321) );
  OAI22XL U1900 ( .A0(n1509), .A1(n1793), .B0(n1324), .B1(n1792), .Y(n1510) );
  OAI22X1 U1901 ( .A0(n1473), .A1(n3106), .B0(n1323), .B1(n3109), .Y(n1511) );
  NAND2X1 U1902 ( .A(n696), .B(n695), .Y(n694) );
  OAI22XL U1903 ( .A0(n3452), .A1(n4081), .B0(n3515), .B1(n4082), .Y(n3512) );
  OAI22XL U1904 ( .A0(n3517), .A1(n4077), .B0(n4078), .B1(n3516), .Y(n4083) );
  OAI21XL U1905 ( .A0(n2585), .A1(n2586), .B0(n2584), .Y(n785) );
  NAND2BXL U1906 ( .AN(n2810), .B(n1050), .Y(n1049) );
  INVXL U1907 ( .A(n1050), .Y(n1048) );
  NAND2X1 U1908 ( .A(n868), .B(n1001), .Y(n2957) );
  XOR3X2 U1909 ( .A(n2955), .B(n2954), .C(n2953), .Y(n2965) );
  INVXL U1910 ( .A(n3356), .Y(n2944) );
  NAND2X1 U1911 ( .A(n775), .B(n774), .Y(n2945) );
  NOR2X1 U1912 ( .A(Q[23]), .B(butt_a_real[4]), .Y(n3611) );
  NAND2XL U1913 ( .A(n2917), .B(n2918), .Y(n765) );
  NAND2XL U1914 ( .A(n3366), .B(n3365), .Y(n1108) );
  INVXL U1915 ( .A(n3365), .Y(n1110) );
  OAI22XL U1916 ( .A0(n3263), .A1(n3275), .B0(n3276), .B1(n3273), .Y(n3281) );
  OAI2BB1XL U1917 ( .A0N(n2362), .A1N(n2361), .B0(n1880), .Y(n3563) );
  NAND2XL U1918 ( .A(n3488), .B(n1998), .Y(n1999) );
  OAI21XL U1919 ( .A0(n3488), .A1(n1998), .B0(butt_b_real[17]), .Y(n2000) );
  OAI22XL U1920 ( .A0(n2240), .A1(n4077), .B0(n2270), .B1(n4078), .Y(n2256) );
  OAI22XL U1921 ( .A0(n2242), .A1(n3445), .B0(n2267), .B1(n3446), .Y(n2254) );
  OAI22XL U1922 ( .A0(n2241), .A1(n2361), .B0(n2268), .B1(n2362), .Y(n2255) );
  INVXL U1923 ( .A(n2311), .Y(n2310) );
  NAND2X1 U1924 ( .A(n842), .B(n843), .Y(n841) );
  NAND2XL U1925 ( .A(n2134), .B(n2133), .Y(n1064) );
  NAND2X1 U1926 ( .A(n1027), .B(n1030), .Y(n1026) );
  INVXL U1927 ( .A(n1057), .Y(n722) );
  OAI2BB1X2 U1928 ( .A0N(n1057), .A1N(n779), .B0(n2047), .Y(n1056) );
  OAI22XL U1929 ( .A0(n1411), .A1(n3271), .B0(n1416), .B1(n3269), .Y(n1421) );
  NAND2X1 U1930 ( .A(n781), .B(n780), .Y(n1568) );
  NAND2XL U1931 ( .A(n782), .B(n1486), .Y(n780) );
  OAI21X1 U1932 ( .A0(n1486), .A1(n782), .B0(n1485), .Y(n781) );
  OR2XL U1933 ( .A(n2656), .B(n2655), .Y(n2659) );
  NOR2X1 U1934 ( .A(n3496), .B(n3497), .Y(n3484) );
  NAND2XL U1935 ( .A(Q[30]), .B(butt_a_real[11]), .Y(n4389) );
  NAND2XL U1936 ( .A(Q[29]), .B(butt_a_real[10]), .Y(n4384) );
  OAI21XL U1937 ( .A0(n3740), .A1(n3728), .B0(n3727), .Y(n4387) );
  NOR2X1 U1938 ( .A(Q[26]), .B(butt_a_real[7]), .Y(n4337) );
  NAND2XL U1939 ( .A(Q[26]), .B(butt_a_real[7]), .Y(n4338) );
  OAI2BB1X2 U1940 ( .A0N(n2869), .A1N(n2870), .B0(n2805), .Y(n2960) );
  XOR2XL U1941 ( .A(n4336), .B(n3610), .Y(n4404) );
  NOR2X1 U1942 ( .A(Q[24]), .B(butt_a_real[5]), .Y(n3618) );
  NAND2XL U1943 ( .A(Q[24]), .B(butt_a_real[5]), .Y(n3619) );
  NAND2XL U1944 ( .A(Q[23]), .B(butt_a_real[4]), .Y(n3614) );
  XOR2XL U1945 ( .A(n1017), .B(n3516), .Y(n3559) );
  XOR2XL U1946 ( .A(n4053), .B(n3660), .Y(n4187) );
  INVXL U1947 ( .A(cs[1]), .Y(n924) );
  XNOR2XL U1948 ( .A(n2388), .B(n2089), .Y(n4604) );
  XNOR2XL U1949 ( .A(n3699), .B(n3698), .Y(n4603) );
  XNOR2XL U1950 ( .A(n4058), .B(n4057), .Y(n4583) );
  OAI21XL U1951 ( .A0(n4053), .A1(n4052), .B0(n4051), .Y(n4058) );
  XOR2XL U1952 ( .A(n3672), .B(n3671), .Y(n4606) );
  OAI21XL U1953 ( .A0(n4510), .A1(n4509), .B0(n4508), .Y(n4511) );
  XNOR2XL U1954 ( .A(n3501), .B(n3500), .Y(n4434) );
  XNOR2XL U1955 ( .A(n3735), .B(n3734), .Y(n4451) );
  XOR2XL U1956 ( .A(n3740), .B(n3739), .Y(n4366) );
  INVXL U1957 ( .A(n4404), .Y(n4356) );
  XOR2XL U1958 ( .A(n4247), .B(n3948), .Y(n4565) );
  NAND2X1 U1959 ( .A(n1461), .B(n1460), .Y(n4415) );
  INVXL U1960 ( .A(n3528), .Y(n4017) );
  NAND2XL U1961 ( .A(n3565), .B(n3564), .Y(n3569) );
  NAND2XL U1962 ( .A(Q[16]), .B(butt_a_imag[16]), .Y(n2380) );
  INVXL U1963 ( .A(n2371), .Y(n3459) );
  NOR2BX2 U1964 ( .AN(n2339), .B(n2289), .Y(n2291) );
  XOR2XL U1965 ( .A(n2393), .B(n2392), .Y(n4601) );
  AOI21XL U1966 ( .A0(n2388), .A1(n2387), .B0(n2386), .Y(n2393) );
  NAND2XL U1967 ( .A(n3811), .B(n605), .Y(n2070) );
  INVX2 U1968 ( .A(n4671), .Y(n2057) );
  NAND2XL U1969 ( .A(n4667), .B(n4665), .Y(n4666) );
  NAND2XL U1970 ( .A(in_out_cnt[8]), .B(n4663), .Y(n4660) );
  NAND2XL U1971 ( .A(n3806), .B(n838), .Y(n3847) );
  INVXL U1972 ( .A(n1011), .Y(n838) );
  AND2XL U1973 ( .A(is_row), .B(n3803), .Y(n3795) );
  BUFX1 U1974 ( .A(n924), .Y(n3965) );
  OAI22XL U1975 ( .A0(n3782), .A1(n3781), .B0(n3780), .B1(n3779), .Y(n3783) );
  XOR2XL U1976 ( .A(IN_VALID), .B(n3778), .Y(n3782) );
  OAI2BB2XL U1977 ( .B0(n3810), .B1(n3821), .A0N(n3786), .A1N(n4666), .Y(n3807) );
  NAND2XL U1978 ( .A(n3779), .B(n3811), .Y(n2101) );
  NAND2XL U1979 ( .A(n4040), .B(n4039), .Y(n4041) );
  INVXL U1980 ( .A(n4038), .Y(n4040) );
  AOI211XL U1981 ( .A0(n4602), .A1(n4496), .B0(n4495), .C0(n4494), .Y(n4497)
         );
  AOI21XL U1982 ( .A0(n4467), .A1(n3465), .B0(n3464), .Y(n3466) );
  NAND2XL U1983 ( .A(n3723), .B(n3722), .Y(n3724) );
  NAND2XL U1984 ( .A(n4331), .B(n4330), .Y(n4332) );
  INVXL U1985 ( .A(n4329), .Y(n4331) );
  NAND2XL U1986 ( .A(n3601), .B(n3600), .Y(n3602) );
  INVXL U1987 ( .A(n721), .Y(n3601) );
  NAND2XL U1988 ( .A(n4310), .B(n4309), .Y(n4311) );
  OAI2BB1XL U1989 ( .A0N(FFT2D_IN_R[3]), .A1N(n4600), .B0(n4315), .Y(n4316) );
  AOI21XL U1990 ( .A0(FFT2D_IN_I[3]), .A1(n4608), .B0(n4314), .Y(n4315) );
  NAND2XL U1991 ( .A(n3596), .B(n3595), .Y(n3597) );
  NAND2XL U1992 ( .A(n3604), .B(n3592), .Y(n3605) );
  OAI2BB1XL U1993 ( .A0N(n4614), .A1N(n3923), .B0(n3922), .Y(n3924) );
  NAND2XL U1994 ( .A(n3899), .B(n3926), .Y(n3927) );
  NAND2XL U1995 ( .A(n3901), .B(n650), .Y(n3903) );
  AOI211XL U1996 ( .A0(n4226), .A1(n4605), .B0(n4225), .C0(n4224), .Y(n4227)
         );
  NOR2X1 U1997 ( .A(n4220), .B(n4552), .Y(n4225) );
  AND2X1 U1998 ( .A(n2330), .B(n2344), .Y(n1115) );
  NAND4XL U1999 ( .A(n4200), .B(n4199), .C(n4198), .D(n4197), .Y(n4201) );
  XOR2XL U2000 ( .A(n3682), .B(n3681), .Y(n3956) );
  NAND2XL U2001 ( .A(n3680), .B(n3679), .Y(n3681) );
  AOI21XL U2002 ( .A0(n4540), .A1(n4538), .B0(n3678), .Y(n3682) );
  INVXL U2003 ( .A(n4537), .Y(n3678) );
  OAI2BB1XL U2004 ( .A0N(n4614), .A1N(n3954), .B0(n3953), .Y(n3955) );
  NAND2XL U2005 ( .A(n3958), .B(n713), .Y(n3959) );
  NAND3XL U2006 ( .A(n4106), .B(lay_cnt[1]), .C(n4644), .Y(n4646) );
  INVXL U2007 ( .A(n3829), .Y(n4624) );
  NAND2XL U2008 ( .A(n4103), .B(n4626), .Y(n4638) );
  NAND2XL U2009 ( .A(n3785), .B(n3811), .Y(n3821) );
  INVXL U2010 ( .A(n3784), .Y(n3785) );
  AOI211XL U2011 ( .A0(n3846), .A1(lay_cnt[4]), .B0(n3819), .C0(n3818), .Y(
        n3828) );
  NAND2XL U2012 ( .A(n4661), .B(in_out_cnt[2]), .Y(n3823) );
  NOR2X1 U2013 ( .A(IN_VALID), .B(n3822), .Y(n4649) );
  NAND2XL U2014 ( .A(n4646), .B(n3834), .Y(n4621) );
  NAND2XL U2015 ( .A(n4106), .B(n3827), .Y(n4626) );
  NAND2XL U2016 ( .A(n4661), .B(in_out_cnt[0]), .Y(n4109) );
  INVXL U2017 ( .A(n1215), .Y(n947) );
  OAI21X1 U2018 ( .A0(n1007), .A1(n1006), .B0(n1334), .Y(n1475) );
  NAND2XL U2019 ( .A(n1336), .B(butt_a_imag[8]), .Y(n1334) );
  INVXL U2020 ( .A(butt_a_imag[7]), .Y(n1006) );
  NAND2XL U2021 ( .A(n1154), .B(n1153), .Y(n1167) );
  XOR2X1 U2022 ( .A(n1475), .B(n808), .Y(n1340) );
  XOR2X1 U2023 ( .A(butt_b_imag[9]), .B(butt_a_imag[9]), .Y(n1476) );
  INVX2 U2024 ( .A(butt_b_imag[8]), .Y(n1336) );
  INVXL U2025 ( .A(butt_b_imag[7]), .Y(n1337) );
  NAND2X2 U2026 ( .A(n999), .B(n998), .Y(n1271) );
  NAND2BX1 U2027 ( .AN(butt_b_imag[6]), .B(butt_a_imag[6]), .Y(n998) );
  OAI21X1 U2028 ( .A0(n1156), .A1(butt_a_imag[6]), .B0(butt_a_imag[5]), .Y(
        n999) );
  INVXL U2029 ( .A(butt_a_real[6]), .Y(n1195) );
  NAND2XL U2030 ( .A(n2431), .B(n2430), .Y(n2461) );
  NAND2XL U2031 ( .A(n2436), .B(butt_a_real[12]), .Y(n2430) );
  OAI21XL U2032 ( .A0(n2436), .A1(butt_a_real[12]), .B0(butt_a_real[11]), .Y(
        n2431) );
  NAND2XL U2033 ( .A(n2741), .B(n2740), .Y(n2896) );
  NAND2XL U2034 ( .A(n2891), .B(butt_a_real[2]), .Y(n2740) );
  OAI21XL U2035 ( .A0(n2891), .A1(butt_a_real[2]), .B0(butt_a_real[1]), .Y(
        n2741) );
  INVXL U2036 ( .A(butt_b_real[3]), .Y(n2745) );
  INVXL U2037 ( .A(n3177), .Y(n677) );
  XNOR2XL U2038 ( .A(n645), .B(n2512), .Y(n3007) );
  INVX2 U2039 ( .A(n2974), .Y(n1107) );
  NAND2BXL U2040 ( .AN(n3270), .B(n2979), .Y(n2980) );
  NAND2BX1 U2041 ( .AN(n3270), .B(n1749), .Y(n1776) );
  NAND2X1 U2042 ( .A(n768), .B(n2197), .Y(n1670) );
  INVXL U2043 ( .A(n3270), .Y(n768) );
  INVX2 U2044 ( .A(butt_b_imag[10]), .Y(n1518) );
  INVXL U2045 ( .A(butt_b_imag[9]), .Y(n1519) );
  NAND2X1 U2046 ( .A(n1033), .B(n1528), .Y(n2162) );
  NAND2XL U2047 ( .A(n2126), .B(n2127), .Y(n1033) );
  NAND2XL U2048 ( .A(n1527), .B(n1526), .Y(n1604) );
  NAND2XL U2049 ( .A(n1529), .B(butt_b_real[10]), .Y(n1526) );
  OAI21XL U2050 ( .A0(n1529), .A1(butt_b_real[10]), .B0(butt_b_real[9]), .Y(
        n1527) );
  INVXL U2051 ( .A(butt_a_real[11]), .Y(n1634) );
  INVXL U2052 ( .A(butt_a_real[12]), .Y(n1633) );
  NAND2XL U2053 ( .A(n1328), .B(n1327), .Y(n1482) );
  NAND2XL U2054 ( .A(n1330), .B(butt_b_real[8]), .Y(n1327) );
  OAI21XL U2055 ( .A0(n1330), .A1(butt_b_real[8]), .B0(butt_b_real[7]), .Y(
        n1328) );
  INVXL U2056 ( .A(butt_a_real[10]), .Y(n1529) );
  INVXL U2057 ( .A(butt_a_real[9]), .Y(n1530) );
  NAND2XL U2058 ( .A(n1631), .B(n1630), .Y(n1699) );
  NAND2XL U2059 ( .A(n1633), .B(butt_b_real[12]), .Y(n1630) );
  OAI21XL U2060 ( .A0(n1633), .A1(butt_b_real[12]), .B0(n681), .Y(n1631) );
  XNOR2X1 U2061 ( .A(butt_a_real[13]), .B(n2466), .Y(n2462) );
  INVXL U2062 ( .A(butt_a_real[14]), .Y(n1750) );
  INVXL U2063 ( .A(butt_a_real[13]), .Y(n1751) );
  XNOR2X2 U2064 ( .A(butt_a_real[14]), .B(butt_b_real[14]), .Y(n2467) );
  INVXL U2065 ( .A(butt_b_imag[11]), .Y(n1657) );
  NAND2X2 U2066 ( .A(n1067), .B(n897), .Y(n961) );
  OAI21X2 U2067 ( .A0(butt_b_imag[2]), .A1(n966), .B0(n965), .Y(n1222) );
  INVXL U2068 ( .A(butt_a_imag[2]), .Y(n966) );
  OAI21X1 U2069 ( .A0(n1165), .A1(butt_a_imag[2]), .B0(n2057), .Y(n965) );
  INVX2 U2070 ( .A(butt_b_imag[2]), .Y(n1165) );
  INVXL U2071 ( .A(n3270), .Y(n673) );
  INVXL U2072 ( .A(n1608), .Y(n634) );
  NAND2XL U2073 ( .A(n582), .B(n2900), .Y(n747) );
  XOR2XL U2074 ( .A(n1013), .B(n3237), .Y(n1577) );
  NAND2XL U2075 ( .A(n1189), .B(n1188), .Y(n1270) );
  NAND2XL U2076 ( .A(n1195), .B(butt_b_real[6]), .Y(n1188) );
  OAI21XL U2077 ( .A0(n1195), .A1(butt_b_real[6]), .B0(butt_b_real[5]), .Y(
        n1189) );
  INVXL U2078 ( .A(butt_a_real[3]), .Y(n1180) );
  INVXL U2079 ( .A(butt_a_real[5]), .Y(n1196) );
  NAND2XL U2080 ( .A(n1179), .B(butt_b_real[4]), .Y(n1171) );
  OAI21X1 U2081 ( .A0(n1179), .A1(butt_b_real[4]), .B0(butt_b_real[3]), .Y(
        n1172) );
  XOR2X2 U2082 ( .A(butt_b_imag[7]), .B(butt_a_imag[7]), .Y(n1272) );
  INVX2 U2083 ( .A(butt_b_imag[6]), .Y(n1156) );
  INVXL U2084 ( .A(butt_b_imag[5]), .Y(n1157) );
  XNOR2X1 U2085 ( .A(n3164), .B(n1528), .Y(n1828) );
  XNOR2X1 U2086 ( .A(n3234), .B(n2830), .Y(n1829) );
  XNOR2X1 U2087 ( .A(n645), .B(n657), .Y(n1773) );
  XNOR2X1 U2088 ( .A(n3451), .B(n2979), .Y(n1757) );
  INVXL U2089 ( .A(n1652), .Y(n1653) );
  INVXL U2090 ( .A(n2264), .Y(n942) );
  XNOR2XL U2091 ( .A(n725), .B(n1528), .Y(n1702) );
  INVXL U2092 ( .A(n1701), .Y(n716) );
  XOR2X1 U2093 ( .A(n627), .B(n573), .Y(n1677) );
  INVXL U2094 ( .A(n2695), .Y(n2696) );
  XNOR2XL U2095 ( .A(n1017), .B(n2757), .Y(n2695) );
  XNOR2XL U2096 ( .A(n755), .B(n2711), .Y(n2712) );
  XOR2XL U2097 ( .A(n1017), .B(n574), .Y(n3447) );
  XOR2X2 U2098 ( .A(n1766), .B(butt_a_imag[14]), .Y(n1768) );
  NAND2XL U2099 ( .A(n1656), .B(butt_a_imag[12]), .Y(n1647) );
  OAI21XL U2100 ( .A0(n1656), .A1(butt_a_imag[12]), .B0(butt_a_imag[11]), .Y(
        n1648) );
  INVXL U2101 ( .A(butt_b_real[15]), .Y(n2452) );
  XNOR2X1 U2102 ( .A(n3451), .B(n2757), .Y(n2664) );
  INVXL U2103 ( .A(n2526), .Y(n2527) );
  OAI2BB1XL U2104 ( .A0N(n2839), .A1N(n2836), .B0(n2830), .Y(n2694) );
  XNOR2XL U2105 ( .A(n2849), .B(n2757), .Y(n2486) );
  OAI2BB1XL U2106 ( .A0N(n3087), .A1N(n3085), .B0(n2475), .Y(n2482) );
  INVXL U2107 ( .A(n2474), .Y(n2475) );
  OAI2BB1XL U2108 ( .A0N(n2940), .A1N(n2938), .B0(n2900), .Y(n2481) );
  XNOR2XL U2109 ( .A(n3014), .B(n2757), .Y(n2497) );
  XOR2X1 U2110 ( .A(n579), .B(n901), .Y(n2498) );
  XNOR2X1 U2111 ( .A(n3270), .B(n4076), .Y(n2415) );
  OAI22XL U2112 ( .A0(n2472), .A1(n3450), .B0(n3449), .B1(n2566), .Y(n2557) );
  NAND2X1 U2113 ( .A(n2619), .B(n1051), .Y(n714) );
  XNOR2XL U2114 ( .A(n949), .B(n2432), .Y(n2571) );
  XNOR2X1 U2115 ( .A(n3054), .B(n2830), .Y(n2564) );
  XNOR2XL U2116 ( .A(n580), .B(n2757), .Y(n2565) );
  XNOR2XL U2117 ( .A(n2783), .B(n657), .Y(n2756) );
  XNOR2X1 U2118 ( .A(n2976), .B(n591), .Y(n2789) );
  NAND2XL U2119 ( .A(n895), .B(n891), .Y(n890) );
  INVXL U2120 ( .A(n2755), .Y(n891) );
  NAND2XL U2121 ( .A(n1097), .B(n583), .Y(n1096) );
  XNOR2X1 U2122 ( .A(n769), .B(n2432), .Y(n2792) );
  XNOR2XL U2123 ( .A(n627), .B(n2900), .Y(n2791) );
  NAND2XL U2124 ( .A(n2420), .B(n2419), .Y(n2510) );
  NAND2XL U2125 ( .A(n2504), .B(butt_a_real[8]), .Y(n2419) );
  OAI21XL U2126 ( .A0(butt_a_real[8]), .A1(n2504), .B0(butt_a_real[7]), .Y(
        n2420) );
  AND2X2 U2127 ( .A(n2501), .B(n2500), .Y(n1069) );
  NAND2XL U2128 ( .A(n2634), .B(butt_a_real[6]), .Y(n2500) );
  NOR2X1 U2129 ( .A(n2505), .B(butt_a_real[7]), .Y(n2499) );
  INVXL U2130 ( .A(butt_b_real[8]), .Y(n2504) );
  INVXL U2131 ( .A(butt_b_real[7]), .Y(n2505) );
  XNOR2X2 U2132 ( .A(n2424), .B(butt_a_real[9]), .Y(n2511) );
  INVXL U2133 ( .A(butt_b_real[6]), .Y(n2634) );
  INVXL U2134 ( .A(butt_b_real[5]), .Y(n2635) );
  INVX2 U2135 ( .A(butt_b_imag[4]), .Y(n1224) );
  INVXL U2136 ( .A(n3085), .Y(n732) );
  NAND2BX1 U2137 ( .AN(n645), .B(n2432), .Y(n2833) );
  XOR2X1 U2138 ( .A(n588), .B(n3004), .Y(n2936) );
  XNOR2X1 U2139 ( .A(n3164), .B(n2979), .Y(n3107) );
  NAND2XL U2140 ( .A(n990), .B(n583), .Y(n988) );
  XNOR2XL U2141 ( .A(n627), .B(n2979), .Y(n3108) );
  XNOR2XL U2142 ( .A(n3270), .B(n3173), .Y(n3178) );
  INVXL U2143 ( .A(butt_b_real[1]), .Y(n2892) );
  XNOR2XL U2144 ( .A(n1038), .B(n3173), .Y(n2994) );
  OAI22XL U2145 ( .A0(n3092), .A1(n3093), .B0(n3091), .B1(n986), .Y(n3128) );
  INVX1 U2146 ( .A(n2989), .Y(n1024) );
  INVXL U2147 ( .A(n996), .Y(n995) );
  XNOR2X1 U2148 ( .A(n578), .B(n3181), .Y(n3090) );
  NAND2XL U2149 ( .A(n1748), .B(n1747), .Y(n1788) );
  NAND2XL U2150 ( .A(n1750), .B(butt_b_real[14]), .Y(n1747) );
  OAI21XL U2151 ( .A0(n1750), .A1(butt_b_real[14]), .B0(butt_b_real[13]), .Y(
        n1748) );
  INVX2 U2152 ( .A(butt_a_real[15]), .Y(n1882) );
  XOR2X2 U2153 ( .A(butt_b_imag[15]), .B(butt_a_imag[15]), .Y(n1770) );
  INVXL U2154 ( .A(butt_b_imag[15]), .Y(n1893) );
  XOR2XL U2155 ( .A(n1017), .B(n901), .Y(n2363) );
  INVXL U2156 ( .A(n2265), .Y(n2266) );
  XNOR2XL U2157 ( .A(n755), .B(n2567), .Y(n2300) );
  XNOR2X1 U2158 ( .A(n3054), .B(n1954), .Y(n1783) );
  XNOR2XL U2159 ( .A(n580), .B(n2900), .Y(n1779) );
  XNOR2X1 U2160 ( .A(n769), .B(n2900), .Y(n1711) );
  XNOR2X1 U2161 ( .A(n3164), .B(n1954), .Y(n1710) );
  XNOR2XL U2162 ( .A(n949), .B(n591), .Y(n1775) );
  XNOR2XL U2163 ( .A(n1036), .B(n1749), .Y(n2233) );
  OAI2BB1XL U2164 ( .A0N(n2199), .A1N(n2198), .B0(n2197), .Y(n2262) );
  XNOR2XL U2165 ( .A(n2976), .B(n1749), .Y(n2203) );
  XNOR2XL U2166 ( .A(n580), .B(n2567), .Y(n2182) );
  OAI22XL U2167 ( .A0(n2181), .A1(n2264), .B0(n2115), .B1(n2263), .Y(n2165) );
  XNOR2X1 U2168 ( .A(n3239), .B(n2567), .Y(n1898) );
  XNOR2XL U2169 ( .A(n3009), .B(n2900), .Y(n1943) );
  OAI22X1 U2170 ( .A0(n1889), .A1(n3110), .B0(n1941), .B1(n3112), .Y(n1936) );
  NAND2X1 U2171 ( .A(n667), .B(n926), .Y(n2163) );
  NAND2XL U2172 ( .A(n2940), .B(n2938), .Y(n926) );
  INVX1 U2173 ( .A(n2162), .Y(n1032) );
  OAI22XL U2174 ( .A0(n2024), .A1(n3558), .B0(n3557), .B1(n3542), .Y(n2107) );
  OAI22X1 U2175 ( .A0(n2025), .A1(n4078), .B0(n4077), .B1(n3516), .Y(n2106) );
  NAND2BX1 U2176 ( .AN(n3270), .B(n3556), .Y(n2024) );
  NAND2X1 U2177 ( .A(n1004), .B(n1003), .Y(n1920) );
  NAND2XL U2178 ( .A(n1005), .B(n944), .Y(n1003) );
  OAI21XL U2179 ( .A0(n1005), .A1(n944), .B0(n1835), .Y(n1004) );
  NOR2BXL U2180 ( .AN(n645), .B(n3446), .Y(n1877) );
  OR2XL U2181 ( .A(n1943), .B(n2938), .Y(n1063) );
  NAND2XL U2182 ( .A(n1062), .B(n582), .Y(n1061) );
  INVXL U2183 ( .A(n2938), .Y(n1060) );
  XNOR2XL U2184 ( .A(n3201), .B(n657), .Y(n1911) );
  XNOR2X1 U2185 ( .A(n3250), .B(n2567), .Y(n1959) );
  XNOR2XL U2186 ( .A(n949), .B(n2830), .Y(n2014) );
  NAND2BXL U2187 ( .AN(n3270), .B(n1173), .Y(n1253) );
  XNOR2XL U2188 ( .A(n645), .B(n3173), .Y(n1256) );
  NAND2XL U2189 ( .A(n1176), .B(n1175), .Y(n1201) );
  NAND2XL U2190 ( .A(n1209), .B(butt_b_real[2]), .Y(n1175) );
  OAI21XL U2191 ( .A0(n1209), .A1(butt_b_real[2]), .B0(butt_b_real[1]), .Y(
        n1176) );
  XOR2XL U2192 ( .A(n1166), .B(n1165), .Y(n1078) );
  XNOR2X2 U2193 ( .A(n1225), .B(butt_a_imag[3]), .Y(n1223) );
  NAND2X1 U2194 ( .A(n796), .B(n793), .Y(n792) );
  INVXL U2195 ( .A(n3269), .Y(n793) );
  INVXL U2196 ( .A(n3275), .Y(n720) );
  INVXL U2197 ( .A(n1094), .Y(n1093) );
  INVXL U2198 ( .A(n3271), .Y(n795) );
  OR2X1 U2199 ( .A(n1279), .B(n3269), .Y(n797) );
  XNOR2X1 U2200 ( .A(n2788), .B(n1606), .Y(n1357) );
  XOR2X1 U2201 ( .A(n1073), .B(n585), .Y(n1322) );
  OAI22XL U2202 ( .A0(n1757), .A1(n3109), .B0(n1762), .B1(n3106), .Y(n1835) );
  INVXL U2203 ( .A(n1718), .Y(n1641) );
  INVXL U2204 ( .A(n1673), .Y(n1713) );
  NOR2X1 U2205 ( .A(n1706), .B(n3112), .Y(n742) );
  XOR2X2 U2206 ( .A(n1756), .B(n941), .Y(n1781) );
  OAI22X1 U2207 ( .A0(n1702), .A1(n2126), .B0(n1782), .B1(n2127), .Y(n1780) );
  INVX1 U2208 ( .A(n1733), .Y(n696) );
  OAI22XL U2209 ( .A0(n1544), .A1(n3109), .B0(n1591), .B1(n3106), .Y(n1588) );
  OAI22X1 U2210 ( .A0(n1610), .A1(n1956), .B0(n1560), .B1(n1955), .Y(n1612) );
  OAI22XL U2211 ( .A0(n1716), .A1(n1793), .B0(n1792), .B1(n1602), .Y(n1667) );
  OAI22X1 U2212 ( .A0(n1679), .A1(n2127), .B0(n2126), .B1(n1601), .Y(n1668) );
  OAI22X1 U2213 ( .A0(n1600), .A1(n3177), .B0(n3179), .B1(n1087), .Y(n1669) );
  NAND2XL U2214 ( .A(n2406), .B(n2405), .Y(n2445) );
  NAND2XL U2215 ( .A(n2451), .B(butt_a_real[16]), .Y(n2405) );
  OAI21XL U2216 ( .A0(n2451), .A1(butt_a_real[16]), .B0(butt_a_real[15]), .Y(
        n2406) );
  XNOR2XL U2217 ( .A(n755), .B(n2674), .Y(n3515) );
  OAI22XL U2218 ( .A0(n2664), .A1(n2763), .B0(n2695), .B1(n2765), .Y(n2693) );
  OAI22XL U2219 ( .A0(n2665), .A1(n2753), .B0(n2755), .B1(n592), .Y(n2692) );
  OAI22XL U2220 ( .A0(n2717), .A1(n4082), .B0(n2701), .B1(n4081), .Y(n2714) );
  OAI22XL U2221 ( .A0(n2698), .A1(n3445), .B0(n2713), .B1(n3446), .Y(n2716) );
  OAI22XL U2222 ( .A0(n2718), .A1(n4078), .B0(n2699), .B1(n4077), .Y(n2715) );
  ADDFX2 U2223 ( .A(n2688), .B(n2687), .CI(n2686), .CO(n2724), .S(n2684) );
  OAI22XL U2224 ( .A0(n2673), .A1(n3445), .B0(n2698), .B1(n3446), .Y(n2687) );
  XNOR2XL U2225 ( .A(n580), .B(n2674), .Y(n2676) );
  ADDFHX1 U2226 ( .A(n2478), .B(n2477), .CI(n2476), .CO(n2545), .S(n2553) );
  OAI22X1 U2227 ( .A0(n2442), .A1(n2846), .B0(n2473), .B1(n2883), .Y(n2478) );
  ADDFX2 U2228 ( .A(n2691), .B(n2690), .CI(n2689), .CO(n2723), .S(n2704) );
  OAI22XL U2229 ( .A0(n2660), .A1(n4077), .B0(n2699), .B1(n4078), .Y(n2691) );
  NAND2X1 U2230 ( .A(n982), .B(n981), .Y(n2666) );
  NAND2XL U2231 ( .A(n2532), .B(n983), .Y(n981) );
  OAI21XL U2232 ( .A0(n2532), .A1(n983), .B0(n2531), .Y(n982) );
  OAI22XL U2233 ( .A0(n2529), .A1(n2753), .B0(n2665), .B1(n2755), .Y(n2671) );
  OAI22X1 U2234 ( .A0(n2673), .A1(n3446), .B0(n900), .B1(n3445), .Y(n2670) );
  OR2X1 U2235 ( .A(n2487), .B(n4077), .Y(n984) );
  OR2XL U2236 ( .A(n2530), .B(n4078), .Y(n985) );
  OAI22XL U2237 ( .A0(n2486), .A1(n2763), .B0(n2528), .B1(n2765), .Y(n2532) );
  INVXL U2238 ( .A(n2550), .Y(n1105) );
  INVXL U2239 ( .A(n2955), .Y(n800) );
  OAI22X1 U2240 ( .A0(n2401), .A1(n4078), .B0(n4077), .B1(n3516), .Y(n2496) );
  NAND2BXL U2241 ( .AN(n3270), .B(n4076), .Y(n2401) );
  XOR2X2 U2242 ( .A(n2554), .B(n699), .Y(n2589) );
  NOR2BX1 U2243 ( .AN(n645), .B(n4082), .Y(n2577) );
  OAI22XL U2244 ( .A0(n2580), .A1(n3085), .B0(n2514), .B1(n3087), .Y(n2575) );
  NAND2XL U2245 ( .A(n2628), .B(n2627), .Y(n2629) );
  OAI21XL U2246 ( .A0(n2628), .A1(n2627), .B0(n2626), .Y(n2630) );
  OAI22XL U2247 ( .A0(n2770), .A1(n3085), .B0(n2580), .B1(n3087), .Y(n2645) );
  NAND2X1 U2248 ( .A(n701), .B(n700), .Y(n2647) );
  OR2X1 U2249 ( .A(n2614), .B(n2615), .Y(n2644) );
  INVXL U2250 ( .A(n2771), .Y(n684) );
  OAI22XL U2251 ( .A0(n2735), .A1(n2846), .B0(n2617), .B1(n2883), .Y(n2626) );
  NAND2X2 U2252 ( .A(n896), .B(n893), .Y(n2627) );
  OAI22XL U2253 ( .A0(n2595), .A1(n2765), .B0(n2766), .B1(n2763), .Y(n2620) );
  OAI22XL U2254 ( .A0(n2769), .A1(n3087), .B0(n2828), .B1(n3085), .Y(n2786) );
  OAI22XL U2255 ( .A0(n2738), .A1(n2839), .B0(n2784), .B1(n2836), .Y(n2785) );
  NAND2X1 U2256 ( .A(n776), .B(n3338), .Y(n774) );
  OAI22X1 U2257 ( .A0(n2829), .A1(n2883), .B0(n2848), .B1(n2846), .Y(n2856) );
  NAND2XL U2258 ( .A(n3346), .B(n2906), .Y(n2912) );
  INVXL U2259 ( .A(n2918), .Y(n767) );
  OAI22X1 U2260 ( .A0(n2862), .A1(n3110), .B0(n2827), .B1(n3112), .Y(n2878) );
  XOR2X1 U2261 ( .A(n949), .B(n973), .Y(n2930) );
  XNOR2X1 U2262 ( .A(n2937), .B(n3173), .Y(n2929) );
  OAI22XL U2263 ( .A0(n2915), .A1(n3109), .B0(n2905), .B1(n3106), .Y(n3347) );
  OAI22XL U2264 ( .A0(n3165), .A1(n3269), .B0(n2987), .B1(n3271), .Y(n2995) );
  OAI22XL U2265 ( .A0(n3013), .A1(n3091), .B0(n3012), .B1(n3092), .Y(n3020) );
  OAI22XL U2266 ( .A0(n3202), .A1(n3259), .B0(n3167), .B1(n3261), .Y(n3204) );
  OAI22XL U2267 ( .A0(n3200), .A1(n3254), .B0(n3168), .B1(n3256), .Y(n3203) );
  OAI22XL U2268 ( .A0(n3168), .A1(n3254), .B0(n3023), .B1(n3256), .Y(n3171) );
  XNOR2XL U2269 ( .A(n769), .B(n3258), .Y(n3202) );
  NAND2BXL U2270 ( .AN(n3239), .B(n2974), .Y(n3268) );
  NAND2BXL U2271 ( .AN(n3265), .B(n594), .Y(n3266) );
  XOR2XL U2272 ( .A(n1073), .B(n575), .Y(n3236) );
  XNOR2XL U2273 ( .A(n580), .B(n2974), .Y(n3235) );
  XNOR2XL U2274 ( .A(n3234), .B(n2974), .Y(n3264) );
  XNOR2XL U2275 ( .A(n745), .B(n594), .Y(n3272) );
  XNOR2XL U2276 ( .A(n3250), .B(n2974), .Y(n3276) );
  XNOR2XL U2277 ( .A(n3201), .B(n2974), .Y(n3263) );
  INVXL U2278 ( .A(n688), .Y(n686) );
  OAI22XL U2279 ( .A0(n3106), .A1(n3059), .B0(n2967), .B1(n3109), .Y(n3060) );
  OAI22XL U2280 ( .A0(n3177), .A1(n3067), .B0(n3066), .B1(n3179), .Y(n3136) );
  INVX2 U2281 ( .A(butt_b_imag[16]), .Y(n1892) );
  INVXL U2282 ( .A(butt_a_real[16]), .Y(n1881) );
  XNOR2XL U2283 ( .A(n3054), .B(n1880), .Y(n2241) );
  XNOR2XL U2284 ( .A(n2976), .B(n1880), .Y(n2268) );
  XOR2XL U2285 ( .A(n773), .B(n901), .Y(n2267) );
  XNOR2XL U2286 ( .A(n3014), .B(n4076), .Y(n2270) );
  XNOR2XL U2287 ( .A(n3164), .B(n3556), .Y(n2269) );
  XOR2XL U2288 ( .A(n1073), .B(n3542), .Y(n2228) );
  NAND2X1 U2289 ( .A(n864), .B(n863), .Y(n1949) );
  NAND2XL U2290 ( .A(n1903), .B(n1904), .Y(n863) );
  OAI21XL U2291 ( .A0(n1903), .A1(n1904), .B0(n865), .Y(n864) );
  OAI22XL U2292 ( .A0(n1958), .A1(n2264), .B0(n1905), .B1(n2263), .Y(n1976) );
  XOR2X2 U2293 ( .A(n1960), .B(n919), .Y(n1975) );
  INVXL U2294 ( .A(n1925), .Y(n842) );
  INVX1 U2295 ( .A(n843), .Y(n840) );
  NAND2XL U2296 ( .A(n1848), .B(n1849), .Y(n789) );
  NAND2BXL U2297 ( .AN(n1823), .B(n1821), .Y(n1826) );
  INVXL U2298 ( .A(n827), .Y(n825) );
  OAI22XL U2299 ( .A0(n2242), .A1(n3446), .B0(n2214), .B1(n3445), .Y(n2245) );
  OAI22XL U2300 ( .A0(n3446), .A1(n2118), .B0(n2029), .B1(n3445), .Y(n2119) );
  OAI22XL U2301 ( .A0(n2027), .A1(n2263), .B0(n2115), .B1(n2264), .Y(n2121) );
  OAI22XL U2302 ( .A0(n1291), .A1(n3273), .B0(n1290), .B1(n3275), .Y(n1298) );
  OAI22X1 U2303 ( .A0(n1289), .A1(n3106), .B0(n1288), .B1(n3109), .Y(n1299) );
  OAI22XL U2304 ( .A0(n1245), .A1(n1607), .B0(n1236), .B1(n1608), .Y(n1248) );
  OAI22XL U2305 ( .A0(n3254), .A1(n1244), .B0(n1237), .B1(n3256), .Y(n1247) );
  OAI22XL U2306 ( .A0(n1297), .A1(n1701), .B0(n1296), .B1(n1700), .Y(n1307) );
  OAI22XL U2307 ( .A0(n1312), .A1(n1607), .B0(n1245), .B1(n1608), .Y(n1313) );
  OAI22XL U2308 ( .A0(n1291), .A1(n3275), .B0(n1257), .B1(n3273), .Y(n1315) );
  NAND2BXL U2309 ( .AN(n3239), .B(n594), .Y(n1414) );
  NAND2BXL U2310 ( .AN(n3265), .B(n1243), .Y(n1413) );
  XOR2XL U2311 ( .A(n1074), .B(n1076), .Y(n1394) );
  XNOR2XL U2312 ( .A(n3234), .B(n594), .Y(n1412) );
  XNOR2XL U2313 ( .A(n745), .B(n1243), .Y(n1415) );
  XNOR2XL U2314 ( .A(n3250), .B(n594), .Y(n1416) );
  XNOR2XL U2315 ( .A(n3201), .B(n594), .Y(n1411) );
  OAI22XL U2316 ( .A0(n1263), .A1(n3269), .B0(n1279), .B1(n3271), .Y(n1303) );
  OAI22XL U2317 ( .A0(n1295), .A1(n3177), .B0(n1264), .B1(n3179), .Y(n1302) );
  OAI22XL U2318 ( .A0(n1593), .A1(n3112), .B0(n1517), .B1(n3110), .Y(n1595) );
  OAI22XL U2319 ( .A0(n1516), .A1(n1700), .B0(n1592), .B1(n1701), .Y(n1596) );
  NAND2XL U2320 ( .A(n853), .B(n656), .Y(n850) );
  NAND2BXL U2321 ( .AN(n656), .B(n852), .Y(n851) );
  OAI22XL U2322 ( .A0(n2718), .A1(n4077), .B0(n3441), .B1(n4078), .Y(n3439) );
  OAI22XL U2323 ( .A0(n2717), .A1(n4081), .B0(n3452), .B1(n4082), .Y(n3440) );
  OAI22XL U2324 ( .A0(n3441), .A1(n4077), .B0(n3517), .B1(n4078), .Y(n3520) );
  OAI22XL U2325 ( .A0(n2491), .A1(n3449), .B0(n2539), .B1(n3450), .Y(n2536) );
  OAI22X1 U2326 ( .A0(n2489), .A1(n3445), .B0(n3446), .B1(n900), .Y(n2538) );
  NOR2X1 U2327 ( .A(n3729), .B(n4388), .Y(n3482) );
  XOR3X2 U2328 ( .A(n2609), .B(n2610), .C(n2608), .Y(n1002) );
  OAI21XL U2329 ( .A0(n3606), .A1(n3480), .B0(n3479), .Y(n3494) );
  NOR2X1 U2330 ( .A(n4335), .B(n4337), .Y(n3478) );
  NAND2XL U2331 ( .A(n613), .B(n3372), .Y(n3354) );
  NAND2X1 U2332 ( .A(n937), .B(n3373), .Y(n1021) );
  NAND2XL U2333 ( .A(n2840), .B(n2841), .Y(n2924) );
  NAND2XL U2334 ( .A(n2903), .B(n2904), .Y(n2840) );
  OAI21XL U2335 ( .A0(n2903), .A1(n2904), .B0(n2902), .Y(n2841) );
  NAND2XL U2336 ( .A(n3384), .B(n3383), .Y(n3385) );
  NAND2BXL U2337 ( .AN(n3384), .B(n3382), .Y(n3386) );
  OAI21XL U2338 ( .A0(n3910), .A1(n3913), .B0(n3911), .Y(n3915) );
  OAI22XL U2339 ( .A0(n3172), .A1(n3275), .B0(n3199), .B1(n3273), .Y(n3224) );
  OAI22XL U2340 ( .A0(n1263), .A1(n3271), .B0(n3269), .B1(n1310), .Y(n1383) );
  OAI22XL U2341 ( .A0(n3218), .A1(n3256), .B0(n3257), .B1(n3254), .Y(n3299) );
  OAI22XL U2342 ( .A0(n3217), .A1(n3261), .B0(n3262), .B1(n3259), .Y(n3300) );
  OAI22XL U2343 ( .A0(n3264), .A1(n3275), .B0(n3263), .B1(n3273), .Y(n3296) );
  OAI22XL U2344 ( .A0(n3257), .A1(n3256), .B0(n3255), .B1(n3254), .Y(n3298) );
  OAI22X1 U2345 ( .A0(n3262), .A1(n3261), .B0(n3260), .B1(n3259), .Y(n3297) );
  XNOR2XL U2346 ( .A(n725), .B(n594), .Y(n3244) );
  OAI22XL U2347 ( .A0(n3240), .A1(n3261), .B0(n3259), .B1(n588), .Y(n3246) );
  NAND2BXL U2348 ( .AN(n3270), .B(n3253), .Y(n3238) );
  XOR2XL U2349 ( .A(n1038), .B(n575), .Y(n3252) );
  ADDFHX1 U2350 ( .A(n3154), .B(n3153), .CI(n3152), .CO(n3387), .S(n3157) );
  NAND2X1 U2351 ( .A(n3037), .B(n3036), .Y(n3117) );
  NAND2XL U2352 ( .A(n3035), .B(n3034), .Y(n3036) );
  XNOR2XL U2353 ( .A(n755), .B(n4076), .Y(n3541) );
  OAI21X1 U2354 ( .A0(n1015), .A1(n1016), .B0(n1891), .Y(n1939) );
  NAND2XL U2355 ( .A(n1892), .B(butt_a_imag[16]), .Y(n1891) );
  INVXL U2356 ( .A(butt_a_imag[15]), .Y(n1015) );
  XOR2X1 U2357 ( .A(butt_b_imag[17]), .B(butt_a_imag[17]), .Y(n1940) );
  INVXL U2358 ( .A(butt_b_imag[17]), .Y(n2009) );
  XOR2X1 U2359 ( .A(n3530), .B(butt_b_imag[18]), .Y(n2010) );
  NAND2XL U2360 ( .A(n1879), .B(n1878), .Y(n1951) );
  NAND2XL U2361 ( .A(n1881), .B(butt_b_real[16]), .Y(n1878) );
  OAI21XL U2362 ( .A0(n1881), .A1(butt_b_real[16]), .B0(butt_b_real[15]), .Y(
        n1879) );
  INVXL U2363 ( .A(butt_a_real[17]), .Y(n2001) );
  OAI22XL U2364 ( .A0(n2306), .A1(n3557), .B0(n2356), .B1(n3558), .Y(n2354) );
  OAI22XL U2365 ( .A0(n2305), .A1(n4077), .B0(n2365), .B1(n4078), .Y(n2355) );
  OAI22XL U2366 ( .A0(n2356), .A1(n3557), .B0(n3543), .B1(n3558), .Y(n3546) );
  NOR2X1 U2367 ( .A(n2088), .B(n2389), .Y(n2065) );
  OAI21XL U2368 ( .A0(n3656), .A1(n2063), .B0(n2062), .Y(n2083) );
  NOR2X1 U2369 ( .A(n4052), .B(n4054), .Y(n2061) );
  NOR2X1 U2370 ( .A(n3700), .B(n3695), .Y(n2084) );
  OAI22XL U2371 ( .A0(n1393), .A1(n3269), .B0(n1310), .B1(n3271), .Y(n1392) );
  OAI22XL U2372 ( .A0(n1311), .A1(n3256), .B0(n1376), .B1(n3254), .Y(n1391) );
  OAI22XL U2373 ( .A0(n1376), .A1(n3256), .B0(n1410), .B1(n3254), .Y(n1439) );
  XOR2XL U2374 ( .A(n1038), .B(n1076), .Y(n1406) );
  NAND2BXL U2375 ( .AN(n3270), .B(n1606), .Y(n1395) );
  NAND2XL U2376 ( .A(n671), .B(n670), .Y(n1599) );
  NAND2XL U2377 ( .A(n1554), .B(n1555), .Y(n670) );
  NAND2XL U2378 ( .A(Q[10]), .B(butt_a_imag[10]), .Y(n2385) );
  NAND2XL U2379 ( .A(Q[9]), .B(butt_a_imag[9]), .Y(n3696) );
  AOI21XL U2380 ( .A0(n3667), .A1(n3658), .B0(n3657), .Y(n4053) );
  NAND2XL U2381 ( .A(Q[7]), .B(butt_a_imag[7]), .Y(n4055) );
  XNOR3X2 U2382 ( .A(n1057), .B(n2048), .C(n2047), .Y(n2051) );
  OAI2BB1X2 U2383 ( .A0N(n1853), .A1N(n1854), .B0(n1852), .Y(n1859) );
  NAND2XL U2384 ( .A(Q[8]), .B(butt_a_imag[8]), .Y(n3701) );
  NOR2X1 U2385 ( .A(Q[8]), .B(butt_a_imag[8]), .Y(n3700) );
  NAND2XL U2386 ( .A(Q[1]), .B(n2057), .Y(n3942) );
  NAND2XL U2387 ( .A(Q[5]), .B(butt_a_imag[5]), .Y(n3669) );
  NAND2XL U2388 ( .A(Q[4]), .B(butt_a_imag[4]), .Y(n3664) );
  ADDFXL U2389 ( .A(n4517), .B(n4516), .CI(n4515), .CO(n4519), .S(n4086) );
  INVXL U2390 ( .A(n4518), .Y(n4517) );
  OAI2BB1XL U2391 ( .A0N(n4082), .A1N(n4081), .B0(n4080), .Y(n4516) );
  AOI21XL U2392 ( .A0(n3981), .A1(n3979), .B0(n3485), .Y(n4450) );
  NOR2XL U2393 ( .A(n4463), .B(n4459), .Y(n4466) );
  OR2XL U2394 ( .A(Q[33]), .B(butt_a_real[14]), .Y(n3979) );
  NAND2XL U2395 ( .A(Q[32]), .B(butt_a_real[13]), .Y(n3983) );
  NAND2XL U2396 ( .A(n2599), .B(n2600), .Y(n2524) );
  NAND2XL U2397 ( .A(Q[31]), .B(butt_a_real[12]), .Y(n3498) );
  NAND2XL U2398 ( .A(Q[3]), .B(butt_a_imag[3]), .Y(n4249) );
  OAI2BB1X2 U2399 ( .A0N(n2957), .A1N(n1102), .B0(n2651), .Y(n2963) );
  NAND2XL U2400 ( .A(n2958), .B(n2956), .Y(n2651) );
  OR2XL U2401 ( .A(n2956), .B(n2958), .Y(n1102) );
  NAND2XL U2402 ( .A(n2965), .B(n649), .Y(n738) );
  NAND2XL U2403 ( .A(n884), .B(n883), .Y(n649) );
  NAND2XL U2404 ( .A(Q[28]), .B(butt_a_real[9]), .Y(n3732) );
  OAI21XL U2405 ( .A0(n2944), .A1(n2943), .B0(n2942), .Y(n3375) );
  INVXL U2406 ( .A(n3357), .Y(n2943) );
  NAND2XL U2407 ( .A(Q[27]), .B(butt_a_real[8]), .Y(n3737) );
  NAND2XL U2408 ( .A(Q[20]), .B(butt_a_real[1]), .Y(n3911) );
  NAND2XL U2409 ( .A(Q[22]), .B(butt_a_real[3]), .Y(n4278) );
  NAND2XL U2410 ( .A(Q[21]), .B(butt_a_real[2]), .Y(n4274) );
  NAND2XL U2411 ( .A(Q[2]), .B(butt_a_imag[2]), .Y(n4245) );
  NOR2XL U2412 ( .A(Q[2]), .B(butt_a_imag[2]), .Y(n4246) );
  NOR2X1 U2413 ( .A(n3292), .B(n3291), .Y(n3295) );
  AOI21XL U2414 ( .A0(n3279), .A1(n3290), .B0(n3289), .Y(n3294) );
  AND2XL U2415 ( .A(n3288), .B(n3287), .Y(n3289) );
  OAI2BB1XL U2416 ( .A0N(n2315), .A1N(n2314), .B0(n2313), .Y(n2350) );
  NAND2BXL U2417 ( .AN(n2312), .B(n2310), .Y(n2315) );
  INVXL U2418 ( .A(n2339), .Y(n820) );
  NAND2XL U2419 ( .A(n1930), .B(n1931), .Y(n786) );
  NAND2BXL U2420 ( .AN(n1930), .B(n788), .Y(n787) );
  NAND2XL U2421 ( .A(Q[14]), .B(butt_a_imag[14]), .Y(n2074) );
  NAND2XL U2422 ( .A(Q[13]), .B(butt_a_imag[13]), .Y(n4009) );
  NAND2XL U2423 ( .A(n2154), .B(n2153), .Y(n2155) );
  NAND2XL U2424 ( .A(Q[12]), .B(butt_a_imag[12]), .Y(n4047) );
  XNOR3X2 U2425 ( .A(n2139), .B(n2153), .C(n2156), .Y(n2148) );
  NAND2XL U2426 ( .A(Q[11]), .B(butt_a_imag[11]), .Y(n2390) );
  NOR2X1 U2427 ( .A(n1431), .B(n1430), .Y(n1434) );
  AOI21XL U2428 ( .A0(n1419), .A1(n1429), .B0(n1428), .Y(n1433) );
  OR2XL U2429 ( .A(n1427), .B(n1426), .Y(n1429) );
  BUFX1 U2430 ( .A(cs[0]), .Y(n3778) );
  INVXL U2431 ( .A(n3688), .Y(n3690) );
  AND2X2 U2432 ( .A(n4037), .B(n4036), .Y(n647) );
  OAI21X1 U2433 ( .A0(n4034), .A1(n4033), .B0(n4032), .Y(n4035) );
  INVXL U2434 ( .A(n4583), .Y(n4564) );
  BUFX1 U2435 ( .A(n3648), .Y(n4031) );
  NOR2X1 U2436 ( .A(n4418), .B(n4416), .Y(n1465) );
  OAI21X1 U2437 ( .A0(n4418), .A1(n4415), .B0(n4419), .Y(n1464) );
  INVXL U2438 ( .A(n4507), .Y(n4513) );
  NAND2XL U2439 ( .A(n4087), .B(n4086), .Y(n4508) );
  AOI21X1 U2440 ( .A0(n4072), .A1(n3521), .B0(n4071), .Y(n4510) );
  NAND2XL U2441 ( .A(n4068), .B(n3521), .Y(n4506) );
  NAND2XL U2442 ( .A(n3523), .B(n3522), .Y(n4070) );
  NAND2XL U2443 ( .A(Q[35]), .B(butt_a_real[16]), .Y(n3490) );
  INVX2 U2444 ( .A(n3430), .Y(n702) );
  NAND2X1 U2445 ( .A(n3427), .B(n3428), .Y(n4471) );
  INVX2 U2446 ( .A(n3427), .Y(n703) );
  NAND2XL U2447 ( .A(n4466), .B(n4460), .Y(n4461) );
  AOI21X1 U2448 ( .A0(n4467), .A1(n4466), .B0(n4465), .Y(n4468) );
  OAI21XL U2449 ( .A0(n4464), .A1(n4463), .B0(n4462), .Y(n4465) );
  INVXL U2450 ( .A(n4463), .Y(n3972) );
  NAND2XL U2451 ( .A(n3426), .B(n3425), .Y(n4462) );
  AOI21X1 U2452 ( .A0(n4467), .A1(n3969), .B0(n3968), .Y(n3970) );
  AOI21X1 U2453 ( .A0(n571), .A1(n4467), .B0(n3974), .Y(n3975) );
  INVXL U2454 ( .A(n3474), .Y(n3974) );
  XOR2XL U2455 ( .A(n4392), .B(n4391), .Y(n4493) );
  AOI21XL U2456 ( .A0(n4387), .A1(n4386), .B0(n4385), .Y(n4392) );
  INVXL U2457 ( .A(n992), .Y(n4375) );
  NAND2XL U2458 ( .A(n4376), .B(n3717), .Y(n4378) );
  XNOR2XL U2459 ( .A(n4387), .B(n3730), .Y(n4479) );
  INVXL U2460 ( .A(n3719), .Y(n4376) );
  XNOR2XL U2461 ( .A(n4341), .B(n4340), .Y(n4435) );
  OAI21XL U2462 ( .A0(n4336), .A1(n4335), .B0(n4334), .Y(n4341) );
  OAI21XL U2463 ( .A0(n4325), .A1(n721), .B0(n3600), .Y(n4326) );
  BUFX1 U2464 ( .A(n3712), .Y(n3722) );
  INVXL U2465 ( .A(n4435), .Y(n4352) );
  XOR2XL U2466 ( .A(n3622), .B(n3621), .Y(n4393) );
  NAND2X2 U2467 ( .A(n3409), .B(n3408), .Y(n3595) );
  INVXL U2468 ( .A(n3591), .Y(n3604) );
  NAND2X1 U2469 ( .A(n3336), .B(n3335), .Y(n4266) );
  NAND2X1 U2470 ( .A(n1627), .B(n1628), .Y(n4238) );
  NAND2XL U2471 ( .A(n3329), .B(n3328), .Y(n710) );
  OR2X2 U2472 ( .A(n3329), .B(n3328), .Y(n3630) );
  ADDFXL U2473 ( .A(n3576), .B(n3575), .CI(n3574), .CO(n3578), .S(n3564) );
  INVXL U2474 ( .A(n3577), .Y(n3576) );
  OAI2BB1XL U2475 ( .A0N(n4078), .A1N(n4077), .B0(n3560), .Y(n3575) );
  OAI2BB1XL U2476 ( .A0N(n3558), .A1N(n3557), .B0(n3556), .Y(n3577) );
  INVXL U2477 ( .A(n3572), .Y(n3573) );
  OAI21XL U2478 ( .A0(n3571), .A1(n3570), .B0(n3569), .Y(n3572) );
  INVXL U2479 ( .A(n4007), .Y(n4220) );
  NAND2XL U2480 ( .A(n3550), .B(n3549), .Y(n3584) );
  OAI21XL U2481 ( .A0(n2320), .A1(n2289), .B0(n2288), .Y(n2290) );
  INVX2 U2482 ( .A(n2283), .Y(n719) );
  INVX2 U2483 ( .A(n2284), .Y(n718) );
  NOR2X2 U2484 ( .A(n1987), .B(n1986), .Y(n3692) );
  NAND2XL U2485 ( .A(n3998), .B(n4028), .Y(n4002) );
  OAI2BB1X1 U2486 ( .A0N(mode_val), .A1N(n2082), .B0(n4668), .Y(n4608) );
  NOR2X1 U2487 ( .A(n2098), .B(n2332), .Y(n4602) );
  NAND2XL U2488 ( .A(n2372), .B(n2374), .Y(n2376) );
  OAI22XL U2489 ( .A0(n3778), .A1(n3965), .B0(n4644), .B1(n3811), .Y(n2073) );
  INVX2 U2490 ( .A(n3932), .Y(n3958) );
  BUFXL U2491 ( .A(n3957), .Y(n713) );
  NAND2XL U2492 ( .A(n3779), .B(n2100), .Y(n3784) );
  BUFXL U2493 ( .A(n2099), .Y(n2100) );
  NAND2XL U2494 ( .A(n3811), .B(n3965), .Y(n3816) );
  BUFXL U2495 ( .A(n3851), .Y(n672) );
  INVXL U2496 ( .A(Q[0]), .Y(n3867) );
  NAND2XL U2497 ( .A(n604), .B(n3778), .Y(n3637) );
  NAND2BXL U2498 ( .AN(n4669), .B(MODE), .Y(n4668) );
  NAND3XL U2499 ( .A(in_out_cnt[2]), .B(in_out_cnt[1]), .C(in_out_cnt[0]), .Y(
        n3777) );
  NOR2X1 U2500 ( .A(n3849), .B(n3777), .Y(n4656) );
  AOI21XL U2501 ( .A0(n4615), .A1(n4614), .B0(n4613), .Y(n4616) );
  NAND4XL U2502 ( .A(n4612), .B(n4611), .C(n4610), .D(n4609), .Y(n4613) );
  OAI211XL U2503 ( .A0(n4587), .A1(n4586), .B0(n4585), .C0(n4584), .Y(n4588)
         );
  OAI211XL U2504 ( .A0(n4569), .A1(n4568), .B0(n4567), .C0(n4566), .Y(n4570)
         );
  AOI22XL U2505 ( .A0(n4607), .A1(n4565), .B0(n2071), .B1(n4580), .Y(n4566) );
  OAI211XL U2506 ( .A0(n4569), .A1(n4563), .B0(n4555), .C0(n4554), .Y(n4556)
         );
  AOI22XL U2507 ( .A0(n4598), .A1(n4589), .B0(n4572), .B1(n4594), .Y(n4562) );
  AND2XL U2508 ( .A(n4608), .B(FFT2D_IN_R[4]), .Y(n3676) );
  NAND2XL U2509 ( .A(n3956), .B(n4614), .Y(n3683) );
  NAND2XL U2510 ( .A(n4538), .B(n4537), .Y(n4539) );
  OAI2BB1XL U2511 ( .A0N(FFT2D_IN_I[3]), .A1N(n4600), .B0(n4545), .Y(n4546) );
  AOI21XL U2512 ( .A0(FFT2D_IN_R[3]), .A1(n4608), .B0(n4544), .Y(n4545) );
  OAI2BB1XL U2513 ( .A0N(n4530), .A1N(n4529), .B0(n4528), .Y(n4531) );
  NAND2X1 U2514 ( .A(n4523), .B(n4598), .Y(n4534) );
  OAI21X1 U2515 ( .A0(n4514), .A1(n4513), .B0(n4512), .Y(n4522) );
  AOI21X1 U2516 ( .A0(n886), .A1(n4614), .B0(n4096), .Y(n4099) );
  OAI2BB1XL U2517 ( .A0N(n4529), .A1N(n2071), .B0(n4095), .Y(n4096) );
  AOI211XL U2518 ( .A0(n4602), .A1(n4498), .B0(n4094), .C0(n4093), .Y(n4095)
         );
  AOI211XL U2519 ( .A0(n4498), .A1(n4605), .B0(n3505), .C0(n3504), .Y(n3506)
         );
  NAND2XL U2520 ( .A(n4491), .B(n4598), .Y(n4488) );
  AND2X1 U2521 ( .A(n3972), .B(n4462), .Y(n1116) );
  NAND2XL U2522 ( .A(n4460), .B(n3969), .Y(n3971) );
  AOI21XL U2523 ( .A0(n4458), .A1(n4614), .B0(n4457), .Y(n4478) );
  NAND4XL U2524 ( .A(n4456), .B(n4455), .C(n4454), .D(n4453), .Y(n4457) );
  NAND4XL U2525 ( .A(n3990), .B(n3989), .C(n3988), .D(n3987), .Y(n3991) );
  NAND2XL U2526 ( .A(n3654), .B(n3640), .Y(n3655) );
  XNOR2XL U2527 ( .A(n4422), .B(n4421), .Y(n4428) );
  OAI211XL U2528 ( .A0(n4356), .A1(n4568), .B0(n4355), .C0(n4354), .Y(n4357)
         );
  AOI22XL U2529 ( .A0(n4607), .A1(n4353), .B0(n2071), .B1(n4366), .Y(n4354) );
  AOI22XL U2530 ( .A0(n4598), .A1(n4364), .B0(n4441), .B1(n4594), .Y(n4363) );
  AOI22XL U2531 ( .A0(n4598), .A1(n4441), .B0(n4410), .B1(n4594), .Y(n4351) );
  AND2XL U2532 ( .A(n4608), .B(FFT2D_IN_I[4]), .Y(n3626) );
  NAND2XL U2533 ( .A(n3925), .B(n4614), .Y(n3633) );
  OAI2BB2X1 U2534 ( .B0(n4669), .B1(MODE), .A0N(n2082), .A1N(n3858), .Y(n4600)
         );
  XNOR2XL U2535 ( .A(n4298), .B(n4297), .Y(n4304) );
  XOR2XL U2536 ( .A(n4273), .B(n4293), .Y(n4287) );
  XOR2XL U2537 ( .A(n4244), .B(n4417), .Y(n4258) );
  OAI2BB1XL U2538 ( .A0N(n4530), .A1N(n4017), .B0(n3533), .Y(n3534) );
  XOR2X1 U2539 ( .A(n912), .B(n660), .Y(n4019) );
  AND2XL U2540 ( .A(n3548), .B(n3582), .Y(n660) );
  AOI211XL U2541 ( .A0(n4602), .A1(n4206), .B0(n2396), .C0(n2395), .Y(n2397)
         );
  ADDFXL U2542 ( .A(Q[17]), .B(butt_a_imag[17]), .CI(n3527), .CO(n3529), .S(
        n4226) );
  INVXL U2543 ( .A(n2384), .Y(n3527) );
  AOI21XL U2544 ( .A0(n2383), .A1(n2382), .B0(n2381), .Y(n2384) );
  NAND2X1 U2545 ( .A(n4019), .B(n3459), .Y(n4233) );
  AOI21X1 U2546 ( .A0(n4597), .A1(n4614), .B0(n4213), .Y(n4218) );
  NAND4XL U2547 ( .A(n4212), .B(n4211), .C(n4210), .D(n4209), .Y(n4213) );
  AOI21XL U2548 ( .A0(n4589), .A1(n4614), .B0(n4063), .Y(n4064) );
  NAND4XL U2549 ( .A(n4062), .B(n4061), .C(n4060), .D(n4059), .Y(n4063) );
  AOI21XL U2550 ( .A0(n4572), .A1(n4614), .B0(n4192), .Y(n4193) );
  NAND4XL U2551 ( .A(n4191), .B(n4190), .C(n4189), .D(n4188), .Y(n4192) );
  INVXL U2552 ( .A(Q[2]), .Y(n3895) );
  INVX2 U2553 ( .A(n635), .Y(FFT2D_OUT_I[14]) );
  INVX2 U2554 ( .A(n642), .Y(FFT2D_OUT_I[15]) );
  INVX2 U2555 ( .A(n646), .Y(FFT2D_OUT_I[16]) );
  INVX2 U2556 ( .A(n652), .Y(FFT2D_OUT_I[17]) );
  NOR2X1 U2557 ( .A(n3866), .B(n4652), .Y(FFT2D_OUT_I[18]) );
  OAI2BB2X2 U2558 ( .B0(n3866), .B1(n3894), .A0N(Q[1]), .A1N(n570), .Y(
        FFT2D_OUT_R[1]) );
  OAI2BB2X2 U2559 ( .B0(n3866), .B1(n3896), .A0N(Q[2]), .A1N(n570), .Y(
        FFT2D_OUT_R[2]) );
  OAI2BB2X2 U2560 ( .B0(n3866), .B1(n3870), .A0N(Q[5]), .A1N(n570), .Y(
        FFT2D_OUT_R[5]) );
  OAI2BB2X2 U2561 ( .B0(n3866), .B1(n3872), .A0N(Q[6]), .A1N(n570), .Y(
        FFT2D_OUT_R[6]) );
  INVXL U2562 ( .A(n3889), .Y(n641) );
  INVXL U2563 ( .A(n3885), .Y(n651) );
  OAI2BB2X2 U2564 ( .B0(n3866), .B1(n3880), .A0N(Q[13]), .A1N(n570), .Y(
        FFT2D_OUT_R[13]) );
  NOR2XL U2565 ( .A(n4653), .B(n3866), .Y(FFT2D_OUT_R[18]) );
  OAI2BB1XL U2566 ( .A0N(butt_b_imag[1]), .A1N(n4186), .B0(n4183), .Y(n504) );
  OAI2BB1XL U2567 ( .A0N(butt_b_real[15]), .A1N(n4186), .B0(n4151), .Y(n536)
         );
  OAI2BB1XL U2568 ( .A0N(butt_b_imag[15]), .A1N(n4186), .B0(n4169), .Y(n494)
         );
  OAI2BB1XL U2569 ( .A0N(butt_a_real[13]), .A1N(n4147), .B0(n4132), .Y(n531)
         );
  OAI2BB1XL U2570 ( .A0N(n2057), .A1N(n4147), .B0(n1125), .Y(n1126) );
  OAI2BB1XL U2571 ( .A0N(n3488), .A1N(n4147), .B0(n1127), .Y(n1128) );
  OAI2BB1XL U2572 ( .A0N(butt_b_real[0]), .A1N(n4186), .B0(n1129), .Y(n1130)
         );
  OAI2BB1XL U2573 ( .A0N(butt_a_real[9]), .A1N(n4147), .B0(n4136), .Y(n521) );
  OAI2BB1XL U2574 ( .A0N(butt_b_real[2]), .A1N(n4186), .B0(n4164), .Y(n508) );
  OAI2BB1XL U2575 ( .A0N(butt_b_imag[7]), .A1N(n4186), .B0(n4177), .Y(n552) );
  OAI2BB1XL U2576 ( .A0N(butt_b_imag[17]), .A1N(n4186), .B0(n4167), .Y(n498)
         );
  OAI2BB1XL U2577 ( .A0N(butt_a_real[7]), .A1N(n4147), .B0(n4138), .Y(n517) );
  OAI2BB1XL U2578 ( .A0N(butt_a_real[3]), .A1N(n4147), .B0(n4142), .Y(n509) );
  OAI2BB1XL U2579 ( .A0N(butt_a_imag[17]), .A1N(n4147), .B0(n4113), .Y(n497)
         );
  OAI2BB1XL U2580 ( .A0N(butt_a_imag[7]), .A1N(n4147), .B0(n4123), .Y(n551) );
  OAI2BB1XL U2581 ( .A0N(butt_a_imag[0]), .A1N(n4147), .B0(n4127), .Y(n481) );
  OAI2BB1XL U2582 ( .A0N(butt_b_imag[0]), .A1N(n4186), .B0(n4185), .Y(n482) );
  OAI2BB1XL U2583 ( .A0N(butt_a_imag[11]), .A1N(n4147), .B0(n4119), .Y(n485)
         );
  OAI2BB1XL U2584 ( .A0N(butt_b_imag[11]), .A1N(n4186), .B0(n4173), .Y(n486)
         );
  OAI2BB1XL U2585 ( .A0N(butt_a_imag[12]), .A1N(n4147), .B0(n4118), .Y(n487)
         );
  OAI2BB1XL U2586 ( .A0N(butt_b_imag[12]), .A1N(n4186), .B0(n4172), .Y(n488)
         );
  OAI2BB1XL U2587 ( .A0N(butt_a_imag[16]), .A1N(n4147), .B0(n4114), .Y(n495)
         );
  OAI2BB1XL U2588 ( .A0N(butt_b_imag[16]), .A1N(n4186), .B0(n4168), .Y(n496)
         );
  OAI2BB1XL U2589 ( .A0N(butt_b_imag[18]), .A1N(n4186), .B0(n4166), .Y(n500)
         );
  OAI2BB1XL U2590 ( .A0N(butt_a_real[2]), .A1N(n4147), .B0(n4143), .Y(n507) );
  OAI2BB1XL U2591 ( .A0N(butt_a_real[4]), .A1N(n4147), .B0(n4141), .Y(n511) );
  OAI2BB1XL U2592 ( .A0N(butt_a_real[5]), .A1N(n4147), .B0(n4140), .Y(n513) );
  OAI2BB1XL U2593 ( .A0N(butt_a_real[6]), .A1N(n4147), .B0(n4139), .Y(n515) );
  OAI2BB1XL U2594 ( .A0N(butt_b_real[9]), .A1N(n4186), .B0(n4157), .Y(n522) );
  OAI2BB1XL U2595 ( .A0N(butt_b_imag[2]), .A1N(n4186), .B0(n4182), .Y(n526) );
  OAI2BB1XL U2596 ( .A0N(n681), .A1N(n4186), .B0(n4155), .Y(n528) );
  OAI2BB1XL U2597 ( .A0N(butt_b_real[13]), .A1N(n4186), .B0(n4153), .Y(n532)
         );
  OAI2BB1XL U2598 ( .A0N(butt_a_real[14]), .A1N(n4147), .B0(n4131), .Y(n533)
         );
  OAI2BB1XL U2599 ( .A0N(butt_b_real[18]), .A1N(n4186), .B0(n4148), .Y(n542)
         );
  OAI2BB1XL U2600 ( .A0N(butt_b_imag[3]), .A1N(n4186), .B0(n4181), .Y(n544) );
  OAI2BB1XL U2601 ( .A0N(butt_b_imag[4]), .A1N(n4186), .B0(n4180), .Y(n546) );
  OAI2BB1XL U2602 ( .A0N(butt_b_imag[5]), .A1N(n4186), .B0(n4179), .Y(n548) );
  OAI2BB1XL U2603 ( .A0N(butt_b_imag[6]), .A1N(n4186), .B0(n4178), .Y(n550) );
  OAI2BB1XL U2604 ( .A0N(butt_a_imag[8]), .A1N(n4147), .B0(n4122), .Y(n553) );
  OAI2BB1XL U2605 ( .A0N(butt_b_imag[9]), .A1N(n4186), .B0(n4175), .Y(n556) );
  OAI2BB1XL U2606 ( .A0N(n4669), .A1N(mode_val), .B0(n4668), .Y(n557) );
  AOI2BB1XL U2607 ( .A0N(n4184), .A1N(n4145), .B0(n4102), .Y(N1237) );
  OAI31XL U2608 ( .A0(n3815), .A1(n3795), .A2(n3802), .B0(n3788), .Y(n567) );
  NAND2XL U2609 ( .A(n3787), .B(n604), .Y(n3788) );
  OAI2BB1XL U2610 ( .A0N(rst_n), .A1N(n3807), .B0(n3813), .Y(n3787) );
  AOI211XL U2611 ( .A0(n4647), .A1(n4660), .B0(n4664), .C0(n4667), .Y(N1165)
         );
  AOI2BB1XL U2612 ( .A0N(in_out_cnt[8]), .A1N(n4663), .B0(n4662), .Y(N1164) );
  AOI211XL U2613 ( .A0(n3833), .A1(n4657), .B0(n4664), .C0(n4663), .Y(N1163)
         );
  AOI2BB1XL U2614 ( .A0N(in_out_cnt[6]), .A1N(n4659), .B0(n4658), .Y(N1162) );
  AOI211XL U2615 ( .A0(n3837), .A1(n4654), .B0(n4664), .C0(n4659), .Y(N1161)
         );
  AOI2BB1XL U2616 ( .A0N(in_out_cnt[4]), .A1N(n4656), .B0(n4655), .Y(N1160) );
  NAND2XL U2617 ( .A(n4661), .B(n4654), .Y(n4655) );
  AOI211XL U2618 ( .A0(n3849), .A1(n3777), .B0(n4664), .C0(n4656), .Y(N1159)
         );
  OAI22XL U2619 ( .A0(n3775), .A1(n3823), .B0(n3774), .B1(n4109), .Y(N1158) );
  OAI32XL U2620 ( .A0(n4631), .A1(in_out_cnt[0]), .A2(n4664), .B0(
        in_out_cnt[1]), .B1(n4109), .Y(N1157) );
  OAI22XL U2621 ( .A0(n3815), .A1(n3814), .B0(n3813), .B1(n3812), .Y(n566) );
  NOR2X1 U2622 ( .A(n3807), .B(n3806), .Y(n3808) );
  OAI22XL U2623 ( .A0(n3815), .A1(n3797), .B0(n3813), .B1(n3965), .Y(n565) );
  AOI211XL U2624 ( .A0(n3796), .A1(n3795), .B0(n3794), .C0(n3793), .Y(n3797)
         );
  OAI22XL U2625 ( .A0(n3815), .A1(n3805), .B0(n3813), .B1(n618), .Y(n564) );
  NOR2X1 U2626 ( .A(n3807), .B(n3804), .Y(n3805) );
  AOI21XL U2627 ( .A0(lay_cnt[1]), .A1(n3776), .B0(IN_VALID), .Y(WEN) );
  OAI2BB1X1 U2628 ( .A0N(n4594), .A1N(n4597), .B0(n3711), .Y(D_imag[8]) );
  INVXL U2629 ( .A(n620), .Y(n4593) );
  AOI21XL U2630 ( .A0(n4589), .A1(n4596), .B0(n4588), .Y(n4590) );
  NAND2XL U2631 ( .A(n4597), .B(n4598), .Y(n4591) );
  AOI211XL U2632 ( .A0(n4600), .A1(FFT2D_IN_I[6]), .B0(n4571), .C0(n4570), .Y(
        n4576) );
  NAND2XL U2633 ( .A(n4573), .B(n4614), .Y(n4574) );
  NAND2XL U2634 ( .A(n4572), .B(n4596), .Y(n4575) );
  AOI211XL U2635 ( .A0(n4600), .A1(FFT2D_IN_I[5]), .B0(n4557), .C0(n4556), .Y(
        n4561) );
  NAND2XL U2636 ( .A(n4558), .B(n4614), .Y(n4559) );
  NAND2XL U2637 ( .A(n4615), .B(n4596), .Y(n4560) );
  AOI211XL U2638 ( .A0(n4600), .A1(FFT2D_IN_I[4]), .B0(n3676), .C0(n3675), .Y(
        n3684) );
  OAI211XL U2639 ( .A0(n4551), .A1(n4592), .B0(n4550), .C0(n4549), .Y(
        D_imag[3]) );
  NAND2XL U2640 ( .A(n4615), .B(n4598), .Y(n4549) );
  AOI211XL U2641 ( .A0(n4614), .A1(n4548), .B0(n4547), .C0(n4546), .Y(n4550)
         );
  XNOR2XL U2642 ( .A(n4540), .B(n4539), .Y(n4548) );
  NAND4X1 U2643 ( .A(n4536), .B(n4535), .C(n4533), .D(n4534), .Y(D_real[18])
         );
  NAND2X1 U2644 ( .A(n4505), .B(n4594), .Y(n4535) );
  AOI21X1 U2645 ( .A0(n4532), .A1(n4614), .B0(n4531), .Y(n4533) );
  AOI21XL U2646 ( .A0(n879), .A1(n4614), .B0(n4499), .Y(n4500) );
  AOI22X1 U2647 ( .A0(n4491), .A1(n4594), .B0(n4490), .B1(n4596), .Y(n4501) );
  OAI2BB1XL U2648 ( .A0N(n2071), .A1N(n4498), .B0(n4497), .Y(n4499) );
  NAND4X1 U2649 ( .A(n4489), .B(n4488), .C(n4487), .D(n4486), .Y(D_real[14])
         );
  NAND2XL U2650 ( .A(n4490), .B(n4594), .Y(n4487) );
  AOI21XL U2651 ( .A0(n4485), .A1(n4614), .B0(n4484), .Y(n4489) );
  NAND2XL U2652 ( .A(n4490), .B(n4598), .Y(n4477) );
  NAND2XL U2653 ( .A(n4532), .B(n4594), .Y(n4476) );
  NAND2XL U2654 ( .A(n599), .B(n4596), .Y(n3993) );
  AOI21XL U2655 ( .A0(n4364), .A1(n4614), .B0(n3991), .Y(n3992) );
  NAND2XL U2656 ( .A(n886), .B(n4594), .Y(n3994) );
  NAND2XL U2657 ( .A(n599), .B(n4594), .Y(n4443) );
  NAND2XL U2658 ( .A(n886), .B(n4598), .Y(n4445) );
  AOI211XL U2659 ( .A0(n4573), .A1(n4596), .B0(n4430), .C0(n4429), .Y(n4431)
         );
  OAI2BB1XL U2660 ( .A0N(n4614), .A1N(n4428), .B0(n4427), .Y(n4429) );
  NAND2XL U2661 ( .A(n599), .B(n4598), .Y(n4414) );
  NAND2XL U2662 ( .A(n4485), .B(n4594), .Y(n4403) );
  NAND2XL U2663 ( .A(n4458), .B(n4596), .Y(n4402) );
  OAI211XL U2664 ( .A0(n4374), .A1(n4592), .B0(n4373), .C0(n4372), .Y(
        D_real[7]) );
  NAND2XL U2665 ( .A(n4458), .B(n4598), .Y(n4373) );
  AOI21XL U2666 ( .A0(n4441), .A1(n4596), .B0(n4371), .Y(n4372) );
  NAND4XL U2667 ( .A(n4363), .B(n4362), .C(n4361), .D(n4360), .Y(D_real[6]) );
  AOI211XL U2668 ( .A0(n4600), .A1(FFT2D_IN_R[6]), .B0(n4358), .C0(n4357), .Y(
        n4362) );
  NAND2XL U2669 ( .A(n4359), .B(n4614), .Y(n4360) );
  NAND2XL U2670 ( .A(n4410), .B(n4596), .Y(n4361) );
  NAND4XL U2671 ( .A(n4351), .B(n4350), .C(n4349), .D(n4348), .Y(D_real[5]) );
  AOI211XL U2672 ( .A0(n4600), .A1(FFT2D_IN_R[5]), .B0(n4346), .C0(n4345), .Y(
        n4350) );
  NAND2XL U2673 ( .A(n4347), .B(n4614), .Y(n4348) );
  NAND2XL U2674 ( .A(n4399), .B(n4596), .Y(n4349) );
  AOI21XL U2675 ( .A0(n4598), .A1(n4410), .B0(n3635), .Y(n3636) );
  AOI211XL U2676 ( .A0(n4600), .A1(FFT2D_IN_R[4]), .B0(n3626), .C0(n3625), .Y(
        n3634) );
  NAND2XL U2677 ( .A(n4399), .B(n4598), .Y(n4319) );
  AOI211XL U2678 ( .A0(n4614), .A1(n4318), .B0(n4317), .C0(n4316), .Y(n4320)
         );
  XNOR2XL U2679 ( .A(n614), .B(n4311), .Y(n4318) );
  AOI211XL U2680 ( .A0(n4359), .A1(n4596), .B0(n4306), .C0(n4305), .Y(n4307)
         );
  OAI2BB1XL U2681 ( .A0N(n4614), .A1N(n4304), .B0(n4303), .Y(n4305) );
  AOI211XL U2682 ( .A0(n4347), .A1(n4596), .B0(n4289), .C0(n4288), .Y(n4290)
         );
  OAI2BB1XL U2683 ( .A0N(n4614), .A1N(n4287), .B0(n4286), .Y(n4288) );
  AOI211XL U2684 ( .A0(n4558), .A1(n4596), .B0(n4260), .C0(n4259), .Y(n4261)
         );
  OAI2BB1XL U2685 ( .A0N(n4614), .A1N(n4258), .B0(n4257), .Y(n4259) );
  NAND2XL U2686 ( .A(n4347), .B(n4594), .Y(n3928) );
  AOI21XL U2687 ( .A0(n3925), .A1(n4596), .B0(n3924), .Y(n3929) );
  OAI211X1 U2688 ( .A0(n4233), .A1(n4502), .B0(n2400), .C0(n2399), .Y(
        D_imag[15]) );
  AOI21X1 U2689 ( .A0(n4599), .A1(n4614), .B0(n2398), .Y(n2399) );
  AOI22X1 U2690 ( .A0(n4214), .A1(n4596), .B0(n4230), .B1(n4594), .Y(n2400) );
  OAI2BB1XL U2691 ( .A0N(n2071), .A1N(n4226), .B0(n2397), .Y(n2398) );
  AOI21XL U2692 ( .A0(n4614), .A1(n4578), .B0(n4201), .Y(n4202) );
  NAND2XL U2693 ( .A(n655), .B(n4596), .Y(n4203) );
  NAND2XL U2694 ( .A(n4558), .B(n4594), .Y(n3960) );
  AOI21XL U2695 ( .A0(n3956), .A1(n4596), .B0(n3955), .Y(n3961) );
  AOI2BB1XL U2696 ( .A0N(n4677), .A1N(n4646), .B0(n4645), .Y(n4648) );
  AOI2BB1XL U2697 ( .A0N(n4641), .A1N(n4640), .B0(n4639), .Y(n4642) );
  AOI211XL U2698 ( .A0(n4635), .A1(n4644), .B0(n4634), .C0(n4633), .Y(n4637)
         );
  AOI211XL U2699 ( .A0(n4638), .A1(sequence_cnt[2]), .B0(n3831), .C0(n3830), 
        .Y(n3832) );
  OR2XL U2700 ( .A(n3856), .B(n3840), .Y(n3824) );
  AOI211XL U2701 ( .A0(is_row), .A1(n4630), .B0(n4629), .C0(n4628), .Y(n4632)
         );
  OAI21XL U2702 ( .A0(lay_cnt[1]), .A1(n4650), .B0(n4649), .Y(n4651) );
  AOI2BB2X1 U2703 ( .B0(n653), .B1(n3881), .A0N(n3897), .A1N(n3882), .Y(n635)
         );
  OAI22X1 U2704 ( .A0(n2125), .A1(n2198), .B0(n2164), .B1(n2199), .Y(n2170) );
  CLKINVX2 U2705 ( .A(n2612), .Y(n638) );
  NAND2X2 U2706 ( .A(n1640), .B(n1639), .Y(n640) );
  NAND2X1 U2707 ( .A(n815), .B(n584), .Y(n1640) );
  NAND2X1 U2708 ( .A(n903), .B(n1816), .Y(n904) );
  OAI2BB2X2 U2709 ( .B0(n3866), .B1(n3890), .A0N(n641), .A1N(n570), .Y(
        FFT2D_OUT_R[10]) );
  AOI2BB2X1 U2710 ( .B0(n653), .B1(n3883), .A0N(n3897), .A1N(n3884), .Y(n642)
         );
  INVX2 U2711 ( .A(n1136), .Y(n643) );
  XNOR2XL U2712 ( .A(n1017), .B(n657), .Y(n2265) );
  OAI2BB1X2 U2713 ( .A0N(n2872), .A1N(n2871), .B0(n1066), .Y(n2868) );
  XOR3X2 U2714 ( .A(n2871), .B(n2872), .C(n2873), .Y(n3376) );
  NAND2X1 U2715 ( .A(n3717), .B(n934), .Y(n644) );
  NAND2X1 U2716 ( .A(n934), .B(n3717), .Y(n3470) );
  BUFX12 U2717 ( .A(n2569), .Y(n645) );
  OAI22X1 U2718 ( .A0(n3088), .A1(n3087), .B0(n3086), .B1(n3085), .Y(n3130) );
  OAI22X2 U2719 ( .A0(n2770), .A1(n3087), .B0(n2769), .B1(n3085), .Y(n2799) );
  OAI22X1 U2720 ( .A0(n2514), .A1(n3085), .B0(n2474), .B1(n3087), .Y(n2516) );
  OAI22X1 U2721 ( .A0(n2978), .A1(n3184), .B0(n3182), .B1(n2993), .Y(n2999) );
  XNOR2X1 U2722 ( .A(n3164), .B(n591), .Y(n2862) );
  AOI2BB2X1 U2723 ( .B0(n653), .B1(n3875), .A0N(n3897), .A1N(n3876), .Y(n646)
         );
  INVXL U2724 ( .A(n3346), .Y(n2910) );
  XOR2X4 U2725 ( .A(n4042), .B(n4041), .Y(n4589) );
  XOR2X2 U2726 ( .A(n3720), .B(n648), .Y(n4485) );
  AND2X1 U2727 ( .A(n4376), .B(n992), .Y(n648) );
  NAND2X1 U2728 ( .A(n1063), .B(n1061), .Y(n1992) );
  BUFX8 U2729 ( .A(cs[2]), .Y(n3811) );
  OAI2BB2X2 U2730 ( .B0(n3866), .B1(n3886), .A0N(n651), .A1N(n570), .Y(
        FFT2D_OUT_R[11]) );
  AOI2BB2X1 U2731 ( .B0(n653), .B1(n3887), .A0N(n3897), .A1N(n3888), .Y(n652)
         );
  INVX2 U2732 ( .A(n3428), .Y(n902) );
  OAI21X2 U2733 ( .A0(n3908), .A1(n3905), .B0(n3906), .Y(n4272) );
  AOI21X2 U2734 ( .A0(n3311), .A1(n3312), .B0(n3310), .Y(n3908) );
  NAND2X2 U2735 ( .A(n940), .B(n1012), .Y(n654) );
  XNOR3X2 U2736 ( .A(n735), .B(n1027), .C(n2138), .Y(n2145) );
  XOR2X1 U2737 ( .A(n778), .B(n658), .Y(n655) );
  OAI22X1 U2738 ( .A0(n1959), .A1(n3446), .B0(n1898), .B1(n3445), .Y(n1945) );
  NAND4X1 U2739 ( .A(n4101), .B(n4100), .C(n4099), .D(n4098), .Y(D_real[17])
         );
  ADDFHX4 U2740 ( .A(n3003), .B(n3002), .CI(n3001), .CO(n3048), .S(n3188) );
  XNOR2X1 U2741 ( .A(n1036), .B(n2900), .Y(n2563) );
  INVXL U2742 ( .A(n3594), .Y(n3596) );
  ADDFHX4 U2743 ( .A(n3133), .B(n3132), .CI(n3131), .CO(n3365), .S(n3349) );
  INVX8 U2744 ( .A(n690), .Y(n1238) );
  OAI2BB2X2 U2745 ( .B0(n3876), .B1(n3866), .A0N(n3875), .A1N(n570), .Y(
        FFT2D_OUT_R[16]) );
  NAND2X4 U2746 ( .A(n3261), .B(n2895), .Y(n3259) );
  NAND2X1 U2747 ( .A(n2732), .B(n1002), .Y(n1001) );
  NAND2X1 U2748 ( .A(n829), .B(n4598), .Y(n4231) );
  XOR2X1 U2749 ( .A(n736), .B(n1997), .Y(n667) );
  ADDFHX1 U2750 ( .A(n3205), .B(n3204), .CI(n3203), .CO(n3208), .S(n3225) );
  OAI21X2 U2751 ( .A0(n4294), .A1(n4291), .B0(n4295), .Y(n3325) );
  OAI21X4 U2752 ( .A0(n2377), .A1(n2276), .B0(n2378), .Y(n1055) );
  XOR2X4 U2753 ( .A(n1205), .B(n1204), .Y(n1608) );
  OAI2BB1X2 U2754 ( .A0N(n4470), .A1N(n4469), .B0(n4468), .Y(n4474) );
  OAI2BB1X2 U2755 ( .A0N(n666), .A1N(n4469), .B0(n3975), .Y(n783) );
  OAI2BB1X1 U2756 ( .A0N(n751), .A1N(n4469), .B0(n3466), .Y(n711) );
  XNOR2X1 U2757 ( .A(n2885), .B(n1203), .Y(n1205) );
  NAND4X1 U2758 ( .A(n2334), .B(n2335), .C(n2336), .D(n2333), .Y(D_imag[14])
         );
  AOI21X1 U2759 ( .A0(n4595), .A1(n4614), .B0(n2105), .Y(n2336) );
  XOR2X4 U2760 ( .A(n2054), .B(n665), .Y(n4595) );
  OAI2BB2X2 U2761 ( .B0(n3866), .B1(n3865), .A0N(Q[12]), .A1N(n570), .Y(
        FFT2D_OUT_R[12]) );
  OAI2BB2X2 U2762 ( .B0(n3866), .B1(n3863), .A0N(Q[4]), .A1N(n570), .Y(
        FFT2D_OUT_R[4]) );
  OAI2BB2X2 U2763 ( .B0(n3866), .B1(n3888), .A0N(Q[17]), .A1N(n570), .Y(
        FFT2D_OUT_R[17]) );
  OAI2BB2X2 U2764 ( .B0(n3866), .B1(n3884), .A0N(Q[15]), .A1N(n570), .Y(
        FFT2D_OUT_R[15]) );
  OAI2BB2X2 U2765 ( .B0(n3866), .B1(n3882), .A0N(Q[14]), .A1N(n570), .Y(
        FFT2D_OUT_R[14]) );
  OAI2BB2X2 U2766 ( .B0(n3866), .B1(n3874), .A0N(Q[7]), .A1N(n570), .Y(
        FFT2D_OUT_R[7]) );
  XNOR2X4 U2767 ( .A(n1765), .B(n1770), .Y(n657) );
  INVXL U2768 ( .A(n1243), .Y(n1076) );
  NAND2BX2 U2769 ( .AN(n3331), .B(n855), .Y(n3926) );
  INVX2 U2770 ( .A(n591), .Y(n1041) );
  AND2X1 U2771 ( .A(n571), .B(n3474), .Y(n659) );
  INVXL U2772 ( .A(n1606), .Y(n1539) );
  INVX2 U2773 ( .A(n4673), .Y(n3488) );
  INVXL U2774 ( .A(lay_cnt[2]), .Y(n1131) );
  NAND2X2 U2775 ( .A(n3418), .B(n3417), .Y(n992) );
  INVX1 U2776 ( .A(n2757), .Y(n977) );
  INVX1 U2777 ( .A(n2512), .Y(n975) );
  INVX2 U2778 ( .A(n2432), .Y(n976) );
  INVX2 U2779 ( .A(n2979), .Y(n669) );
  NAND2X1 U2780 ( .A(n759), .B(n758), .Y(n2285) );
  INVX2 U2781 ( .A(n1749), .Y(n697) );
  AND2X1 U2782 ( .A(n577), .B(n3977), .Y(n661) );
  AND2X1 U2783 ( .A(n2379), .B(n2378), .Y(n662) );
  AND2X1 U2784 ( .A(n3521), .B(n4070), .Y(n663) );
  XNOR2X2 U2785 ( .A(n1939), .B(n1940), .Y(n2567) );
  INVX2 U2786 ( .A(n2567), .Y(n901) );
  NOR2X2 U2787 ( .A(n1868), .B(n1869), .Y(n3649) );
  AND2X1 U2788 ( .A(n3715), .B(n3714), .Y(n664) );
  AND2X1 U2789 ( .A(n2374), .B(n2276), .Y(n665) );
  BUFX8 U2790 ( .A(n3058), .Y(n1073) );
  XOR2X1 U2791 ( .A(n1209), .B(butt_b_real[2]), .Y(n2885) );
  NOR2X1 U2792 ( .A(n3324), .B(n3323), .Y(n4294) );
  NOR2X2 U2793 ( .A(n3721), .B(n3713), .Y(n3717) );
  INVX2 U2794 ( .A(lay_cnt[3]), .Y(n1138) );
  AND2X1 U2795 ( .A(n4460), .B(n571), .Y(n666) );
  INVX2 U2796 ( .A(n2632), .Y(n979) );
  XNOR3X2 U2797 ( .A(n1603), .B(n2438), .C(n1605), .Y(n2199) );
  NOR2X2 U2798 ( .A(n2371), .B(n2090), .Y(n4614) );
  INVX2 U2799 ( .A(n3516), .Y(n4076) );
  INVX4 U2800 ( .A(Q[37]), .Y(n4653) );
  OAI22X2 U2801 ( .A0(n3200), .A1(n3256), .B0(n3218), .B1(n3254), .Y(n3232) );
  ADDFHX2 U2802 ( .A(n2778), .B(n2777), .CI(n2776), .CO(n2793), .S(n2851) );
  ADDFHX2 U2803 ( .A(n2859), .B(n2858), .CI(n2857), .CO(n2867), .S(n3344) );
  ADDFHX2 U2804 ( .A(n3407), .B(n3406), .CI(n3405), .CO(n3410), .S(n3396) );
  INVX4 U2805 ( .A(n1238), .Y(n726) );
  XNOR2X1 U2806 ( .A(n3270), .B(n657), .Y(n2754) );
  INVX8 U2807 ( .A(n1013), .Y(n3004) );
  XOR2X1 U2808 ( .A(n1252), .B(n1013), .Y(n1479) );
  NAND2X4 U2809 ( .A(n1354), .B(n832), .Y(n1013) );
  OAI22X2 U2810 ( .A0(n2791), .A1(n2938), .B0(n2790), .B1(n2940), .Y(n2797) );
  NOR2X2 U2811 ( .A(n3418), .B(n3417), .Y(n3719) );
  XOR2X1 U2812 ( .A(n3251), .B(n669), .Y(n2983) );
  BUFX8 U2813 ( .A(n3009), .Y(n971) );
  NAND2X4 U2814 ( .A(n3901), .B(n3926), .Y(n4263) );
  XOR3X2 U2815 ( .A(n1555), .B(n1554), .C(n1553), .Y(n1550) );
  BUFX8 U2816 ( .A(n3009), .Y(n972) );
  OAI2BB2X2 U2817 ( .B0(n1355), .B1(n3273), .A0N(n1243), .A1N(n720), .Y(n1489)
         );
  OAI21X4 U2818 ( .A0(n4025), .A1(n2347), .B0(n1052), .Y(n691) );
  NAND2X4 U2819 ( .A(n1054), .B(n2339), .Y(n2347) );
  XOR3X2 U2820 ( .A(n3360), .B(n3358), .C(n3359), .Y(n3407) );
  NAND2XL U2821 ( .A(n1724), .B(n1725), .Y(n674) );
  OAI21X1 U2822 ( .A0(n1724), .A1(n1725), .B0(n1723), .Y(n675) );
  XOR3X2 U2823 ( .A(n1725), .B(n1724), .C(n1723), .Y(n1734) );
  INVX1 U2824 ( .A(n1044), .Y(n676) );
  NAND4X4 U2825 ( .A(n678), .B(n924), .C(n4625), .D(n3811), .Y(n822) );
  NAND2X4 U2826 ( .A(n3750), .B(n3779), .Y(n3817) );
  XNOR2X1 U2827 ( .A(n3201), .B(n3181), .Y(n2993) );
  OAI22X1 U2828 ( .A0(n1955), .A1(n1505), .B0(n1560), .B1(n1956), .Y(n1546) );
  ADDFHX1 U2829 ( .A(n1383), .B(n1382), .CI(n1381), .CO(n1316), .S(n1388) );
  NAND2X4 U2830 ( .A(n3599), .B(n968), .Y(n756) );
  NOR2X4 U2831 ( .A(n4324), .B(n4329), .Y(n968) );
  NAND2X2 U2832 ( .A(n899), .B(n3571), .Y(n898) );
  OAI21X1 U2833 ( .A0(n1848), .A1(n1849), .B0(n1122), .Y(n790) );
  NAND2X2 U2834 ( .A(n3381), .B(n3380), .Y(n3412) );
  ADDFHX4 U2835 ( .A(n1798), .B(n1797), .CI(n1796), .CO(n1901), .S(n1845) );
  XNOR2X1 U2836 ( .A(n1036), .B(n2830), .Y(n2479) );
  ADDFHX1 U2837 ( .A(n1914), .B(n1913), .CI(n1912), .CO(n1970), .S(n1923) );
  ADDFHX2 U2838 ( .A(n3212), .B(n3211), .CI(n3210), .CO(n3326), .S(n3324) );
  NOR2X4 U2839 ( .A(n3325), .B(n679), .Y(n3627) );
  NOR2X2 U2840 ( .A(n680), .B(n4294), .Y(n679) );
  XOR2X1 U2841 ( .A(n3164), .B(n585), .Y(n1506) );
  NOR2BX1 U2842 ( .AN(n645), .B(n3091), .Y(n2991) );
  BUFX2 U2843 ( .A(n1817), .Y(n903) );
  OAI22X1 U2844 ( .A0(n2993), .A1(n3184), .B0(n3185), .B1(n3182), .Y(n3197) );
  OR2X2 U2845 ( .A(n1643), .B(n1642), .Y(n1717) );
  XNOR2X2 U2846 ( .A(n1646), .B(n1768), .Y(n1650) );
  OAI2BB1X2 U2847 ( .A0N(n3091), .A1N(n3092), .B0(n2640), .Y(n2771) );
  OAI2BB2X2 U2848 ( .B0(n1084), .B1(n3254), .A0N(n1079), .A1N(n3253), .Y(n3079) );
  OAI22X1 U2849 ( .A0(n2987), .A1(n3269), .B0(n3005), .B1(n3271), .Y(n2988) );
  OAI2BB1X2 U2850 ( .A0N(n687), .A1N(n3021), .B0(n685), .Y(n3065) );
  XNOR3X2 U2851 ( .A(n3022), .B(n688), .C(n3021), .Y(n3162) );
  AOI2BB2X2 U2852 ( .B0(n689), .B1(n1079), .A0N(n3023), .A1N(n3254), .Y(n688)
         );
  OAI22X1 U2853 ( .A0(n1323), .A1(n3106), .B0(n1289), .B1(n3109), .Y(n1361) );
  XOR3X2 U2854 ( .A(n1002), .B(n2731), .C(n2732), .Y(n2961) );
  OAI21X4 U2855 ( .A0(n1259), .A1(n1186), .B0(n1194), .Y(n690) );
  ADDFHX4 U2856 ( .A(n3341), .B(n3340), .CI(n3339), .CO(n3357), .S(n3372) );
  XNOR2X1 U2857 ( .A(n3251), .B(n3556), .Y(n2114) );
  INVX4 U2858 ( .A(n691), .Y(n914) );
  OAI21X2 U2859 ( .A0(n4027), .A1(n3692), .B0(n3687), .Y(n692) );
  OAI22X1 U2860 ( .A0(n2983), .A1(n3106), .B0(n2982), .B1(n3109), .Y(n2997) );
  NAND2X1 U2861 ( .A(n1733), .B(n1734), .Y(n693) );
  INVXL U2862 ( .A(n1734), .Y(n695) );
  XOR3X2 U2863 ( .A(n1734), .B(n1733), .C(n1732), .Y(n1743) );
  XNOR2X1 U2864 ( .A(n3164), .B(n2197), .Y(n1972) );
  AOI21X1 U2865 ( .A0(n1090), .A1(n4614), .B0(n3534), .Y(n3589) );
  OAI22X1 U2866 ( .A0(n1715), .A1(n1792), .B0(n1764), .B1(n1793), .Y(n1805) );
  XOR2X2 U2867 ( .A(n3251), .B(n697), .Y(n1794) );
  ADDFHX4 U2868 ( .A(n3390), .B(n3389), .CI(n3388), .CO(n3371), .S(n3399) );
  INVX8 U2869 ( .A(n698), .Y(n2975) );
  INVX4 U2870 ( .A(n1503), .Y(n698) );
  OAI2BB1X2 U2871 ( .A0N(n2953), .A1N(n799), .B0(n798), .Y(n2652) );
  NAND2X2 U2872 ( .A(n4472), .B(n3469), .Y(n3433) );
  OAI22XL U2873 ( .A0(n2712), .A1(n3450), .B0(n2697), .B1(n3449), .Y(n2719) );
  INVX8 U2874 ( .A(n704), .Y(n1140) );
  NOR2X4 U2875 ( .A(cs[2]), .B(cs[3]), .Y(n704) );
  NAND2X2 U2876 ( .A(n1552), .B(n1551), .Y(n1621) );
  OAI22X1 U2877 ( .A0(n1764), .A1(n1792), .B0(n1793), .B1(n587), .Y(n1838) );
  OAI22X1 U2878 ( .A0(n1507), .A1(n1607), .B0(n1540), .B1(n1608), .Y(n1558) );
  NOR2X4 U2879 ( .A(n3997), .B(n4003), .Y(n2339) );
  ADDFHX4 U2880 ( .A(n1346), .B(n1345), .CI(n1344), .CO(n1485), .S(n1351) );
  XOR2X1 U2881 ( .A(n736), .B(n3028), .Y(n1070) );
  XNOR2X1 U2882 ( .A(n3201), .B(n2979), .Y(n1323) );
  OAI21X1 U2883 ( .A0(n2824), .A1(n2825), .B0(n2823), .Y(n705) );
  NAND2X2 U2884 ( .A(n1162), .B(n1193), .Y(n1280) );
  CLKINVX8 U2885 ( .A(n1199), .Y(n1193) );
  NAND2X4 U2886 ( .A(n2055), .B(n4625), .Y(n1199) );
  NAND2X1 U2887 ( .A(n1870), .B(n1871), .Y(n4039) );
  XOR3X2 U2888 ( .A(n944), .B(n1005), .C(n1835), .Y(n1840) );
  ADDFHX4 U2889 ( .A(n1693), .B(n1692), .CI(n1691), .CO(n1815), .S(n1739) );
  OAI2BB1X2 U2890 ( .A0N(n3158), .A1N(n708), .B0(n707), .Y(n3332) );
  XOR3X2 U2891 ( .A(n3160), .B(n3159), .C(n3158), .Y(n3329) );
  OAI22X1 U2892 ( .A0(n2563), .A1(n2938), .B0(n2940), .B1(n1997), .Y(n2520) );
  OAI22X1 U2893 ( .A0(n3897), .A1(n3868), .B0(n3867), .B1(n3866), .Y(
        FFT2D_OUT_I[0]) );
  NAND2X4 U2894 ( .A(n4653), .B(n3859), .Y(n3897) );
  OAI22XL U2895 ( .A0(n2528), .A1(n2763), .B0(n2664), .B1(n2765), .Y(n2661) );
  BUFX1 U2896 ( .A(n3817), .Y(n712) );
  XNOR2X1 U2897 ( .A(n3251), .B(n1528), .Y(n1601) );
  XOR2X2 U2898 ( .A(n3251), .B(n573), .Y(n1505) );
  XNOR2X1 U2899 ( .A(n3239), .B(n3253), .Y(n1409) );
  OAI22X1 U2900 ( .A0(n3185), .A1(n3184), .B0(n3183), .B1(n3182), .Y(n3220) );
  ADDFHX1 U2901 ( .A(n3000), .B(n2999), .CI(n2998), .CO(n3189), .S(n3193) );
  NAND2X1 U2902 ( .A(n790), .B(n789), .Y(n1926) );
  XOR2X1 U2903 ( .A(n3164), .B(n901), .Y(n900) );
  CLKINVX2 U2904 ( .A(n714), .Y(n2591) );
  NAND2BXL U2905 ( .AN(n3270), .B(n2567), .Y(n2568) );
  NAND2XL U2906 ( .A(n715), .B(n3181), .Y(n3175) );
  INVX2 U2907 ( .A(n3239), .Y(n715) );
  ADDFHX4 U2908 ( .A(n3096), .B(n3095), .CI(n3094), .CO(n3156), .S(n3119) );
  XNOR2X2 U2909 ( .A(n745), .B(n2567), .Y(n2574) );
  OAI22X4 U2910 ( .A0(n2574), .A1(n3445), .B0(n3446), .B1(n1014), .Y(n2588) );
  OAI21X2 U2911 ( .A0(n1214), .A1(n1199), .B0(n1354), .Y(n717) );
  AND2X2 U2912 ( .A(n3309), .B(n3308), .Y(n3310) );
  NAND2XL U2913 ( .A(n875), .B(n874), .Y(n873) );
  XOR2X2 U2914 ( .A(n2886), .B(n2888), .Y(n2974) );
  ADDFHX1 U2915 ( .A(n3247), .B(n3246), .CI(n3245), .CO(n3302), .S(n3306) );
  AOI21X1 U2916 ( .A0(n4000), .A1(n2339), .B0(n2346), .Y(n2328) );
  ADDFHX1 U2917 ( .A(n2124), .B(n2123), .CI(n2122), .CO(n2150), .S(n2138) );
  AOI21X2 U2918 ( .A0(n1086), .A1(n4614), .B0(n4018), .Y(n4022) );
  NAND4X2 U2919 ( .A(n4023), .B(n4021), .C(n4022), .D(n4020), .Y(D_imag[17])
         );
  ADDFHX4 U2920 ( .A(n3350), .B(n3349), .CI(n3348), .CO(n3389), .S(n3367) );
  NAND2X4 U2921 ( .A(n719), .B(n718), .Y(n2330) );
  ADDFHX1 U2922 ( .A(n1380), .B(n1379), .CI(n1378), .CO(n1381), .S(n1397) );
  NOR2X1 U2923 ( .A(n1273), .B(n3818), .Y(n1275) );
  NAND2X1 U2924 ( .A(n724), .B(n723), .Y(n1864) );
  NOR2BX2 U2925 ( .AN(n3270), .B(n2755), .Y(n2782) );
  INVXL U2926 ( .A(n763), .Y(n762) );
  ADDFHX1 U2927 ( .A(n2262), .B(n2261), .CI(n2260), .CO(n2299), .S(n2257) );
  XOR3X2 U2928 ( .A(n3366), .B(n3365), .C(n3364), .Y(n3392) );
  NOR2BX1 U2929 ( .AN(n3239), .B(n3256), .Y(n1404) );
  NOR2X4 U2930 ( .A(n3433), .B(n4463), .Y(n936) );
  OAI21X2 U2931 ( .A0(n3474), .A1(n3976), .B0(n3977), .Y(n3968) );
  NOR2X4 U2932 ( .A(n3423), .B(n3424), .Y(n3976) );
  ADDFHX2 U2933 ( .A(n2553), .B(n2552), .CI(n2551), .CO(n2522), .S(n2606) );
  NOR2X2 U2934 ( .A(n1011), .B(n837), .Y(n836) );
  ADDFHX4 U2935 ( .A(n3402), .B(n3401), .CI(n3400), .CO(n3403), .S(n3335) );
  OAI22X2 U2936 ( .A0(n2833), .A1(n2883), .B0(n2846), .B1(n976), .Y(n2880) );
  ADDHX2 U2937 ( .A(n2880), .B(n2881), .CO(n2855), .S(n2918) );
  INVX2 U2938 ( .A(cs[2]), .Y(n3812) );
  OAI22XL U2939 ( .A0(n1290), .A1(n3273), .B0(n1355), .B1(n3275), .Y(n1344) );
  ADDFHX4 U2940 ( .A(n3051), .B(n3050), .CI(n3049), .CO(n3096), .S(n3047) );
  OAI22X1 U2941 ( .A0(n1357), .A1(n1608), .B0(n1236), .B1(n1607), .Y(n1320) );
  AOI21X4 U2942 ( .A0(n939), .A1(n811), .B0(n938), .Y(n862) );
  NAND2X4 U2943 ( .A(n845), .B(n764), .Y(n1216) );
  NAND2X4 U2944 ( .A(n2279), .B(n2280), .Y(n3999) );
  OAI21X1 U2945 ( .A0(n1744), .A1(n1746), .B0(n1745), .Y(n724) );
  XOR3X4 U2946 ( .A(n1746), .B(n1745), .C(n1744), .Y(n1628) );
  OAI2BB1X2 U2947 ( .A0N(n1956), .A1N(n1955), .B0(n1954), .Y(n1996) );
  INVX1 U2948 ( .A(n3031), .Y(n1058) );
  OAI22XL U2949 ( .A0(n2915), .A1(n3106), .B0(n3107), .B1(n3109), .Y(n3143) );
  XOR2X1 U2950 ( .A(n4241), .B(n4240), .Y(n4587) );
  NAND2X4 U2951 ( .A(n940), .B(n1012), .Y(n811) );
  ADDFHX4 U2952 ( .A(n1676), .B(n1675), .CI(n1674), .CO(n1712), .S(n1687) );
  INVX2 U2953 ( .A(n2935), .Y(n3073) );
  ADDFHX1 U2954 ( .A(n1566), .B(n1565), .CI(n1564), .CO(n1614), .S(n1569) );
  NAND2BXL U2955 ( .AN(n3270), .B(n2830), .Y(n2832) );
  OAI22X1 U2956 ( .A0(n3107), .A1(n3106), .B0(n3109), .B1(n3108), .Y(n3151) );
  OAI21X4 U2957 ( .A0(n4640), .A1(n1099), .B0(n3812), .Y(n1153) );
  BUFX4 U2958 ( .A(n579), .Y(n725) );
  ADDFHX2 U2959 ( .A(n2589), .B(n2588), .CI(n2587), .CO(n2598), .S(n2613) );
  NAND2X4 U2960 ( .A(n726), .B(n772), .Y(n3058) );
  NAND2X2 U2961 ( .A(n3331), .B(n3332), .Y(n3899) );
  NAND2X1 U2962 ( .A(n744), .B(n1100), .Y(n2648) );
  OAI21X2 U2963 ( .A0(n731), .A1(n730), .B0(n729), .Y(n3424) );
  OAI21X1 U2964 ( .A0(n2603), .A1(n2604), .B0(n2602), .Y(n729) );
  INVX2 U2965 ( .A(n2603), .Y(n730) );
  NOR2X2 U2966 ( .A(n616), .B(n3421), .Y(n3473) );
  NOR2X4 U2967 ( .A(n4263), .B(n4265), .Y(n969) );
  NOR2X4 U2968 ( .A(n3335), .B(n3336), .Y(n4265) );
  INVXL U2969 ( .A(n2340), .Y(n2341) );
  ADDFHX1 U2970 ( .A(n2309), .B(n2308), .CI(n2307), .CO(n2353), .S(n2298) );
  ADDFHX1 U2971 ( .A(n2352), .B(n2351), .CI(n2350), .CO(n2370), .S(n2316) );
  NOR2X4 U2972 ( .A(n1193), .B(n1162), .Y(n1259) );
  OAI21X1 U2973 ( .A0(n2951), .A1(n2952), .B0(n885), .Y(n884) );
  OAI22XL U2974 ( .A0(n3244), .A1(n3269), .B0(n3236), .B1(n3271), .Y(n3303) );
  INVX1 U2975 ( .A(n859), .Y(n856) );
  NAND2X4 U2976 ( .A(n1199), .B(n1162), .Y(n1163) );
  BUFX8 U2977 ( .A(n1162), .Y(n1353) );
  INVXL U2978 ( .A(n4461), .Y(n4470) );
  XNOR2X1 U2979 ( .A(n3201), .B(n2674), .Y(n2488) );
  XNOR2X1 U2980 ( .A(n3201), .B(n2711), .Y(n2566) );
  XOR2X1 U2981 ( .A(n2975), .B(n593), .Y(n2913) );
  OAI2BB1X4 U2982 ( .A0N(n667), .A1N(n582), .B0(n1059), .Y(n2109) );
  INVX4 U2983 ( .A(n1625), .Y(n1012) );
  NOR2X4 U2984 ( .A(n2280), .B(n2279), .Y(n3997) );
  AND2X4 U2985 ( .A(n1282), .B(n1193), .Y(n770) );
  XOR2X4 U2986 ( .A(n2422), .B(n2421), .Y(n3087) );
  INVX3 U2987 ( .A(n1285), .Y(n1071) );
  XNOR2X1 U2988 ( .A(n3004), .B(n3084), .Y(n2474) );
  XNOR3X2 U2989 ( .A(n2134), .B(n2133), .C(n2132), .Y(n735) );
  BUFX2 U2990 ( .A(n1013), .Y(n736) );
  BUFX12 U2991 ( .A(n2849), .Y(n949) );
  INVX1 U2992 ( .A(n2752), .Y(n2835) );
  ADDFHX1 U2993 ( .A(n1917), .B(n1916), .CI(n1915), .CO(n1969), .S(n1900) );
  OAI22X2 U2994 ( .A0(n2443), .A1(n4078), .B0(n2415), .B1(n4077), .Y(n2517) );
  XNOR3X2 U2995 ( .A(n2965), .B(n2966), .C(n740), .Y(n3418) );
  OAI21X2 U2996 ( .A0(n2376), .A1(n4027), .B0(n2375), .Y(n737) );
  AND2X2 U2997 ( .A(n645), .B(n805), .Y(n1342) );
  OAI21X2 U2998 ( .A0(n739), .A1(n740), .B0(n738), .Y(n3420) );
  NOR2X1 U2999 ( .A(n2965), .B(n649), .Y(n739) );
  XNOR3X2 U3000 ( .A(n2956), .B(n2958), .C(n2957), .Y(n740) );
  XOR2X4 U3001 ( .A(n2450), .B(n2449), .Y(n3450) );
  XNOR2X1 U3002 ( .A(n578), .B(n3258), .Y(n3015) );
  INVX2 U3003 ( .A(n1274), .Y(n844) );
  ADDFHX1 U3004 ( .A(n2787), .B(n2786), .CI(n2785), .CO(n2824), .S(n2866) );
  XNOR2X1 U3005 ( .A(n3239), .B(n3181), .Y(n3183) );
  OAI21X1 U3006 ( .A0(n2465), .A1(butt_a_real[14]), .B0(butt_a_real[13]), .Y(
        n2448) );
  NAND3X2 U3007 ( .A(n1164), .B(n961), .C(n831), .Y(n1325) );
  BUFX12 U3008 ( .A(n1325), .Y(n3014) );
  OAI22X1 U3009 ( .A0(n2914), .A1(n2940), .B0(n2941), .B1(n2938), .Y(n3144) );
  ADDFHX1 U3010 ( .A(n3148), .B(n3147), .CI(n3146), .CO(n3366), .S(n3352) );
  XOR2X4 U3011 ( .A(n2408), .B(n2407), .Y(n4082) );
  OAI2BB1X2 U3012 ( .A0N(n3179), .A1N(n3177), .B0(n3173), .Y(n2781) );
  NOR2BX1 U3013 ( .AN(n645), .B(n2883), .Y(n2933) );
  INVXL U3014 ( .A(n2293), .Y(n741) );
  OAI2BB1X2 U3015 ( .A0N(n741), .A1N(n2349), .B0(n2292), .Y(n2319) );
  NAND2X1 U3016 ( .A(n771), .B(n3084), .Y(n2934) );
  ADDFHX1 U3017 ( .A(n3437), .B(n3436), .CI(n3435), .CO(n3457), .S(n3429) );
  AOI21X4 U3018 ( .A0(n1054), .A1(n2346), .B0(n1053), .Y(n1052) );
  NOR2X4 U3019 ( .A(n2345), .B(n2338), .Y(n1054) );
  ADDFHX2 U3020 ( .A(n1743), .B(n1742), .CI(n1741), .CO(n1867), .S(n1865) );
  XNOR3X4 U3021 ( .A(n1573), .B(n1658), .C(n1576), .Y(n2839) );
  XNOR2X1 U3022 ( .A(n645), .B(n2674), .Y(n2429) );
  ADDFHX2 U3023 ( .A(n1599), .B(n1598), .CI(n1597), .CO(n1745), .S(n1620) );
  NOR2BX1 U3024 ( .AN(n645), .B(n2940), .Y(n1563) );
  OAI22X2 U3025 ( .A0(n2848), .A1(n2883), .B0(n2847), .B1(n2846), .Y(n2908) );
  XNOR2X2 U3026 ( .A(n1036), .B(n1606), .Y(n1540) );
  BUFX8 U3027 ( .A(n1274), .Y(n764) );
  XOR3X2 U3028 ( .A(n2668), .B(n2666), .C(n2667), .Y(n2682) );
  AOI2BB1X1 U3029 ( .A0N(n1672), .A1N(n3110), .B0(n742), .Y(n1673) );
  OAI22X1 U3030 ( .A0(n1356), .A1(n3110), .B0(n1508), .B1(n3112), .Y(n1488) );
  INVX1 U3031 ( .A(n2954), .Y(n801) );
  NAND2XL U3032 ( .A(n801), .B(n800), .Y(n799) );
  BUFX12 U3033 ( .A(n3010), .Y(n2976) );
  OAI22X1 U3034 ( .A0(n1890), .A1(n1955), .B0(n1956), .B1(n573), .Y(n1946) );
  OAI21X4 U3035 ( .A0(n3999), .A1(n4003), .B0(n4004), .Y(n2346) );
  XOR2X4 U3036 ( .A(n743), .B(n1111), .Y(n829) );
  NAND3X4 U3037 ( .A(n804), .B(n802), .C(n3582), .Y(n743) );
  XNOR2X1 U3038 ( .A(n1036), .B(n2197), .Y(n2164) );
  OR2X4 U3039 ( .A(n1467), .B(n1466), .Y(n4538) );
  ADDFHX1 U3040 ( .A(n1596), .B(n1595), .CI(n1594), .CO(n1726), .S(n1619) );
  ADDFHX1 U3041 ( .A(n3301), .B(n3300), .CI(n3299), .CO(n3242), .S(n3317) );
  OAI21X1 U3042 ( .A0(n2610), .A1(n2609), .B0(n2608), .Y(n744) );
  BUFX4 U3043 ( .A(n1259), .Y(n1234) );
  OR2X2 U3044 ( .A(n3309), .B(n3308), .Y(n3311) );
  NAND2X1 U3045 ( .A(n835), .B(n4598), .Y(n4023) );
  ADDHX1 U3046 ( .A(n1705), .B(n1704), .CO(n1807), .S(n1714) );
  OAI22X2 U3047 ( .A0(n3005), .A1(n3269), .B0(n575), .B1(n3271), .Y(n3041) );
  XNOR2X1 U3048 ( .A(n3234), .B(n2674), .Y(n2540) );
  NOR2X1 U3049 ( .A(n1226), .B(n1227), .Y(n1229) );
  XNOR2X1 U3050 ( .A(n645), .B(n4076), .Y(n2013) );
  OAI2BB1X2 U3051 ( .A0N(n1701), .A1N(n1700), .B0(n1173), .Y(n1756) );
  ADDFHX2 U3052 ( .A(n3157), .B(n3156), .CI(n3155), .CO(n3336), .S(n3333) );
  ADDFHX2 U3053 ( .A(n3045), .B(n3044), .CI(n3043), .CO(n3075), .S(n3050) );
  BUFX8 U3054 ( .A(n3251), .Y(n745) );
  OAI22X1 U3055 ( .A0(n1592), .A1(n1700), .B0(n1654), .B1(n1701), .Y(n1684) );
  NOR2X4 U3056 ( .A(n1866), .B(n1867), .Y(n3642) );
  NAND2X4 U3057 ( .A(n1533), .B(n2127), .Y(n2126) );
  XOR2X4 U3058 ( .A(n1483), .B(n1484), .Y(n2127) );
  XNOR2X1 U3059 ( .A(n2975), .B(n3084), .Y(n2514) );
  XOR2X2 U3060 ( .A(n1094), .B(n929), .Y(n928) );
  OAI22X2 U3061 ( .A0(n1341), .A1(n3112), .B0(n3110), .B1(n1041), .Y(n1094) );
  XNOR2X2 U3062 ( .A(n733), .B(n2446), .Y(n2450) );
  OAI22X1 U3063 ( .A0(n2570), .A1(n3450), .B0(n3449), .B1(n574), .Y(n2619) );
  OAI22XL U3064 ( .A0(n2846), .A1(n2473), .B0(n2883), .B1(n2526), .Y(n2543) );
  OAI22X1 U3065 ( .A0(n2826), .A1(n3109), .B0(n3106), .B1(n669), .Y(n2778) );
  INVXL U3066 ( .A(n3370), .Y(n3373) );
  OAI21X2 U3067 ( .A0(n3721), .A1(n4379), .B0(n3722), .Y(n3716) );
  XOR2X2 U3068 ( .A(n1478), .B(n1477), .Y(n1524) );
  OAI22XL U3069 ( .A0(n1601), .A1(n2127), .B0(n1541), .B1(n2126), .Y(n1582) );
  NAND2X4 U3070 ( .A(n3901), .B(n861), .Y(n4262) );
  OAI22X1 U3071 ( .A0(n3007), .A1(n3068), .B0(n3056), .B1(n3070), .Y(n3040) );
  NAND2X1 U3072 ( .A(n1948), .B(n1949), .Y(n748) );
  XOR3X2 U3073 ( .A(n1949), .B(n1948), .C(n1947), .Y(n1980) );
  NOR2X2 U3074 ( .A(n1462), .B(n1463), .Y(n4418) );
  OAI22X1 U3075 ( .A0(n1799), .A1(n2755), .B0(n1773), .B1(n2753), .Y(n1837) );
  XNOR3X4 U3076 ( .A(n1758), .B(n1894), .C(n1761), .Y(n3446) );
  OAI22X1 U3077 ( .A0(n1782), .A1(n2126), .B0(n1828), .B1(n2127), .Y(n1798) );
  XNOR2X2 U3078 ( .A(n3250), .B(n2757), .Y(n2764) );
  NAND2X4 U3079 ( .A(n750), .B(n1208), .Y(n2783) );
  ADDFHX1 U3080 ( .A(n1558), .B(n1557), .CI(n1556), .CO(n1616), .S(n1554) );
  INVX2 U3081 ( .A(n1187), .Y(n772) );
  OAI22X1 U3082 ( .A0(n2488), .A1(n4082), .B0(n2458), .B1(n4081), .Y(n2485) );
  XOR2X1 U3083 ( .A(n2772), .B(n2771), .Y(n1010) );
  ADDFHX1 U3084 ( .A(n3151), .B(n3150), .CI(n3149), .CO(n3351), .S(n3140) );
  INVXL U3085 ( .A(n3467), .Y(n751) );
  NAND2X1 U3086 ( .A(n754), .B(n753), .Y(n1968) );
  NAND2XL U3087 ( .A(n1919), .B(n1920), .Y(n753) );
  OAI21X1 U3088 ( .A0(n1919), .A1(n1920), .B0(n1918), .Y(n754) );
  XOR3X2 U3089 ( .A(n1920), .B(n1919), .C(n1918), .Y(n1925) );
  NAND2BX2 U3090 ( .AN(n3270), .B(n2900), .Y(n2901) );
  INVX2 U3091 ( .A(n1233), .Y(n1170) );
  OAI22X1 U3092 ( .A0(n2850), .A1(n3092), .B0(n1072), .B1(n3091), .Y(n2842) );
  OAI2BB1X2 U3093 ( .A0N(n1683), .A1N(n851), .B0(n850), .Y(n1692) );
  XOR2X1 U3094 ( .A(n3201), .B(n576), .Y(n3013) );
  INVX2 U3095 ( .A(n1214), .Y(n1233) );
  OAI22X1 U3096 ( .A0(n2487), .A1(n4078), .B0(n2443), .B1(n4077), .Y(n2477) );
  ADDFHX1 U3097 ( .A(n1399), .B(n1398), .CI(n1397), .CO(n1389), .S(n1452) );
  XOR3X4 U3098 ( .A(n1719), .B(n640), .C(n1717), .Y(n1724) );
  OAI21X4 U3099 ( .A0(n3590), .A1(n756), .B0(n932), .Y(n4469) );
  AOI21X4 U3100 ( .A0(n969), .A1(n3898), .B0(n956), .Y(n3590) );
  NAND4X2 U3101 ( .A(n3587), .B(n3589), .C(n3588), .D(n3586), .Y(D_imag[18])
         );
  ADDFHX4 U3102 ( .A(n1902), .B(n1901), .CI(n1900), .CO(n1981), .S(n1924) );
  XNOR3X2 U3103 ( .A(n2247), .B(n757), .C(n2246), .Y(n2222) );
  INVX2 U3104 ( .A(n2248), .Y(n757) );
  OAI21X1 U3105 ( .A0(n2249), .A1(n2250), .B0(n760), .Y(n759) );
  XOR3X4 U3106 ( .A(n1684), .B(n853), .C(n1683), .Y(n1727) );
  INVX2 U3107 ( .A(n1577), .Y(n1578) );
  OAI2BB1X4 U3108 ( .A0N(n3256), .A1N(n3254), .B0(n1578), .Y(n1675) );
  XNOR2X1 U3109 ( .A(n1038), .B(n3556), .Y(n2178) );
  OAI22X1 U3110 ( .A0(n3175), .A1(n3184), .B0(n3182), .B1(n593), .Y(n3176) );
  NOR2X2 U3111 ( .A(n1134), .B(n3851), .Y(n823) );
  OAI22X1 U3112 ( .A0(n2930), .A1(n3092), .B0(n2850), .B1(n3091), .Y(n2907) );
  XOR3X4 U3113 ( .A(n2917), .B(n2918), .C(n2916), .Y(n3362) );
  XNOR2X2 U3114 ( .A(n2425), .B(n1481), .Y(n1484) );
  OAI21X2 U3115 ( .A0(n1991), .A1(n4027), .B0(n1990), .Y(n2054) );
  XNOR2X2 U3116 ( .A(n3251), .B(n4076), .Y(n2443) );
  INVX1 U3117 ( .A(n2599), .Y(n980) );
  ADDFHX2 U3118 ( .A(n2051), .B(n2050), .CI(n2049), .CO(n2053), .S(n1988) );
  ADDFHX1 U3119 ( .A(n2625), .B(n2624), .CI(n2623), .CO(n2650), .S(n2810) );
  INVX4 U3120 ( .A(n821), .Y(n915) );
  XNOR2X1 U3121 ( .A(n1036), .B(n1954), .Y(n1890) );
  XOR3X2 U3122 ( .A(n3338), .B(n776), .C(n3337), .Y(n3378) );
  AOI21X4 U3123 ( .A0(n934), .A1(n1039), .B0(n1101), .Y(n3471) );
  NOR2X4 U3124 ( .A(n3719), .B(n4380), .Y(n934) );
  INVX4 U3125 ( .A(n2099), .Y(n1141) );
  NAND2XL U3126 ( .A(n4097), .B(n4596), .Y(n4098) );
  OAI21X2 U3127 ( .A0(n4027), .A1(n4002), .B0(n4001), .Y(n4006) );
  XOR2X4 U3128 ( .A(n4006), .B(n1114), .Y(n1086) );
  OAI22X2 U3129 ( .A0(n3015), .A1(n3259), .B0(n3053), .B1(n3261), .Y(n3044) );
  ADDFHX4 U3130 ( .A(n3099), .B(n3098), .CI(n3097), .CO(n3139), .S(n3095) );
  AOI21X4 U3131 ( .A0(n777), .A1(n3931), .B0(n1629), .Y(n3638) );
  NOR2X4 U3132 ( .A(n4235), .B(n4237), .Y(n777) );
  NOR2X4 U3133 ( .A(n823), .B(n1258), .Y(n1231) );
  XOR2X1 U3134 ( .A(n778), .B(n658), .Y(n4219) );
  XNOR2X1 U3135 ( .A(n1036), .B(n1243), .Y(n1355) );
  OAI21X2 U3136 ( .A0(n4027), .A1(n2329), .B0(n2328), .Y(n2331) );
  XNOR2X1 U3137 ( .A(n3250), .B(n3237), .Y(n1410) );
  ADDFHX1 U3138 ( .A(n2152), .B(n2151), .CI(n2150), .CO(n2189), .S(n2149) );
  AOI22X2 U3139 ( .A0(n596), .A1(n845), .B0(n1261), .B1(n764), .Y(n1232) );
  NAND2BX2 U3140 ( .AN(n3270), .B(n1528), .Y(n1534) );
  NAND2X1 U3141 ( .A(n1280), .B(n1046), .Y(n1283) );
  ADDFHX4 U3142 ( .A(n2950), .B(n2949), .CI(n2948), .CO(n3416), .S(n3414) );
  ADDFHX1 U3143 ( .A(n1805), .B(n1804), .CI(n1803), .CO(n1823), .S(n1814) );
  XNOR2X1 U3144 ( .A(n1036), .B(n1791), .Y(n1764) );
  XOR2X4 U3145 ( .A(n2743), .B(n2742), .Y(n3184) );
  ADDFHX1 U3146 ( .A(n2170), .B(n2169), .CI(n2168), .CO(n2219), .S(n2185) );
  INVX2 U3147 ( .A(butt_a_imag[10]), .Y(n1035) );
  ADDFHX1 U3148 ( .A(n1318), .B(n1317), .CI(n1316), .CO(n1366), .S(n1368) );
  XOR3X2 U3149 ( .A(n1486), .B(n1485), .C(n782), .Y(n1500) );
  XOR2X4 U3150 ( .A(n928), .B(n1487), .Y(n782) );
  XNOR2X1 U3151 ( .A(n3251), .B(n3173), .Y(n3180) );
  OAI2BB1X4 U3152 ( .A0N(n1820), .A1N(n1855), .B0(n1819), .Y(n1930) );
  ADDFHX1 U3153 ( .A(n3224), .B(n3223), .CI(n3222), .CO(n3206), .S(n3229) );
  ADDFHX1 U3154 ( .A(n3208), .B(n3207), .CI(n3206), .CO(n3191), .S(n3210) );
  NOR2BX2 U3155 ( .AN(n3270), .B(n2127), .Y(n1538) );
  OAI21X2 U3156 ( .A0(n1518), .A1(butt_a_imag[10]), .B0(butt_a_imag[9]), .Y(
        n1034) );
  OAI21X2 U3157 ( .A0(n3600), .A1(n4329), .B0(n4330), .Y(n967) );
  NOR2X4 U3158 ( .A(n2347), .B(n4024), .Y(n2348) );
  ADDFHX4 U3159 ( .A(n2189), .B(n2188), .CI(n2187), .CO(n2281), .S(n2280) );
  XNOR3X2 U3160 ( .A(n2207), .B(n827), .C(n2206), .Y(n2209) );
  XOR2X4 U3161 ( .A(n783), .B(n661), .Y(n886) );
  NOR2X4 U3162 ( .A(n3411), .B(n3412), .Y(n4329) );
  OAI22X1 U3163 ( .A0(n2178), .A1(n3558), .B0(n2114), .B1(n3557), .Y(n2166) );
  ADDFHX4 U3164 ( .A(n2643), .B(n2644), .CI(n2642), .CO(n2610), .S(n2812) );
  OAI22X2 U3165 ( .A0(n2764), .A1(n2765), .B0(n2758), .B1(n2763), .Y(n2777) );
  OAI21X2 U3166 ( .A0(n4379), .A1(n4378), .B0(n4377), .Y(n4383) );
  NAND2X1 U3167 ( .A(n784), .B(n785), .Y(n2581) );
  NAND2XL U3168 ( .A(n2586), .B(n2585), .Y(n784) );
  XOR3X2 U3169 ( .A(n2586), .B(n2585), .C(n2584), .Y(n2955) );
  OAI2BB1X2 U3170 ( .A0N(n787), .A1N(n1929), .B0(n786), .Y(n1986) );
  XNOR3X4 U3171 ( .A(n1930), .B(n788), .C(n1929), .Y(n1870) );
  ADDFHX4 U3172 ( .A(n1739), .B(n1740), .CI(n1738), .CO(n1862), .S(n1741) );
  ADDFHX4 U3173 ( .A(n1863), .B(n1862), .CI(n1861), .CO(n1869), .S(n1866) );
  XOR3X2 U3174 ( .A(n2016), .B(n2017), .C(n2015), .Y(n2047) );
  XOR3X2 U3175 ( .A(n1849), .B(n1848), .C(n1122), .Y(n1860) );
  ADDFHX1 U3176 ( .A(n1546), .B(n1547), .CI(n1545), .CO(n1585), .S(n1555) );
  NAND2X4 U3177 ( .A(n3967), .B(n936), .Y(n935) );
  OAI22X1 U3178 ( .A0(n1670), .A1(n2199), .B0(n2198), .B1(n1075), .Y(n1705) );
  XOR2X2 U3179 ( .A(n3716), .B(n664), .Y(n4458) );
  NAND2BXL U3180 ( .AN(n645), .B(n3028), .Y(n2981) );
  OAI21X1 U3181 ( .A0(n1696), .A1(n1695), .B0(n1694), .Y(n1698) );
  NAND3X2 U3182 ( .A(n2099), .B(n925), .C(lay_cnt[3]), .Y(n970) );
  CLKINVX8 U3183 ( .A(n1099), .Y(n2099) );
  NAND2X4 U3184 ( .A(cs[1]), .B(cs[0]), .Y(n1099) );
  XOR2X1 U3185 ( .A(n645), .B(n2830), .Y(n1664) );
  OAI21X1 U3186 ( .A0(n1479), .A1(n3271), .B0(n792), .Y(n1490) );
  NAND2X1 U3187 ( .A(n796), .B(n795), .Y(n794) );
  XOR2X4 U3188 ( .A(n3451), .B(n594), .Y(n796) );
  NAND2XL U3189 ( .A(n2954), .B(n2955), .Y(n798) );
  NAND2X4 U3190 ( .A(n807), .B(n3112), .Y(n3110) );
  NAND2XL U3191 ( .A(n3933), .B(n654), .Y(n3934) );
  OAI2BB1X4 U3192 ( .A0N(n812), .A1N(n2196), .B0(n2195), .Y(n2223) );
  NAND2X1 U3193 ( .A(n815), .B(n814), .Y(n877) );
  INVXL U3194 ( .A(n2198), .Y(n814) );
  INVX1 U3195 ( .A(n2109), .Y(n818) );
  INVX4 U3196 ( .A(n2330), .Y(n2338) );
  MXI2X2 U3197 ( .A(n845), .B(n1215), .S0(n821), .Y(n917) );
  NAND2X2 U3198 ( .A(n1231), .B(n1285), .Y(n821) );
  NAND2X4 U3199 ( .A(n970), .B(n822), .Y(n1285) );
  NOR2X4 U3200 ( .A(n1133), .B(n1140), .Y(n1258) );
  OAI2BB1X1 U3201 ( .A0N(n2206), .A1N(n826), .B0(n824), .Y(n2234) );
  NAND2XL U3202 ( .A(n825), .B(n2207), .Y(n824) );
  NAND2BXL U3203 ( .AN(n2207), .B(n827), .Y(n826) );
  NAND2X2 U3204 ( .A(n829), .B(n4596), .Y(n3586) );
  NAND2X1 U3205 ( .A(n829), .B(n4594), .Y(n4021) );
  NAND2X4 U3206 ( .A(n830), .B(n1067), .Y(n1207) );
  NAND2X2 U3207 ( .A(n835), .B(n4594), .Y(n3588) );
  XOR2X4 U3208 ( .A(n898), .B(n1112), .Y(n835) );
  INVX4 U3209 ( .A(n836), .Y(n1139) );
  NOR2X2 U3210 ( .A(n1138), .B(cs[1]), .Y(n837) );
  AND2X4 U3211 ( .A(n1786), .B(n1785), .Y(n843) );
  NAND2XL U3212 ( .A(n1831), .B(n848), .Y(n846) );
  OAI21XL U3213 ( .A0(n1831), .A1(n848), .B0(n1830), .Y(n847) );
  XOR3X2 U3214 ( .A(n848), .B(n1831), .C(n1830), .Y(n1846) );
  NOR2X2 U3215 ( .A(cs[1]), .B(cs[3]), .Y(n3752) );
  INVXL U3216 ( .A(n3926), .Y(n3900) );
  NAND2XL U3217 ( .A(n859), .B(n858), .Y(n857) );
  INVXL U3218 ( .A(n3184), .Y(n858) );
  NAND2X2 U3219 ( .A(n3902), .B(n3899), .Y(n861) );
  NAND2X2 U3220 ( .A(n3333), .B(n3334), .Y(n3902) );
  OR2X4 U3221 ( .A(n3333), .B(n3334), .Y(n3901) );
  OAI21X4 U3222 ( .A0(n4262), .A1(n4265), .B0(n4266), .Y(n956) );
  NAND2X4 U3223 ( .A(n3070), .B(n2509), .Y(n3068) );
  OAI21X4 U3224 ( .A0(n862), .A1(n4237), .B0(n4238), .Y(n1629) );
  OAI21XL U3225 ( .A0(n4236), .A1(n4235), .B0(n862), .Y(n4241) );
  AOI2BB2X2 U3226 ( .B0(n867), .B1(n584), .A0N(n1795), .A1N(n2198), .Y(n866)
         );
  INVX1 U3227 ( .A(n1909), .Y(n867) );
  NAND2X4 U3228 ( .A(n870), .B(n1956), .Y(n1955) );
  XNOR3X4 U3229 ( .A(n1269), .B(n2506), .C(n869), .Y(n1956) );
  NAND2XL U3230 ( .A(n1781), .B(n876), .Y(n872) );
  NAND2BX1 U3231 ( .AN(n1778), .B(n584), .Y(n878) );
  NAND2XL U3232 ( .A(n879), .B(n4594), .Y(n4412) );
  NAND2XL U3233 ( .A(n879), .B(n4598), .Y(n4401) );
  NAND2XL U3234 ( .A(n879), .B(n4596), .Y(n4444) );
  NAND2X4 U3235 ( .A(n1080), .B(n882), .Y(n3254) );
  NAND2X2 U3236 ( .A(n884), .B(n883), .Y(n2966) );
  NAND2X1 U3237 ( .A(n2951), .B(n2952), .Y(n883) );
  XOR3X2 U3238 ( .A(n2952), .B(n2951), .C(n885), .Y(n2959) );
  NAND2X1 U3239 ( .A(n1215), .B(n897), .Y(n1206) );
  NAND2X4 U3240 ( .A(n1046), .B(n1274), .Y(n897) );
  OAI21X2 U3241 ( .A0(n1816), .A1(n903), .B0(n1815), .Y(n905) );
  XOR3X2 U3242 ( .A(n1817), .B(n1816), .C(n1815), .Y(n1863) );
  XOR2X4 U3243 ( .A(n910), .B(n908), .Y(n2264) );
  NAND2X2 U3244 ( .A(n1214), .B(n1259), .Y(n916) );
  NAND2X4 U3245 ( .A(n1142), .B(n1276), .Y(n1214) );
  NOR2X4 U3246 ( .A(n3419), .B(n3420), .Y(n4380) );
  NOR2X1 U3247 ( .A(butt_a_imag[15]), .B(n1893), .Y(n1758) );
  NAND2X1 U3248 ( .A(n2274), .B(n2275), .Y(n2378) );
  NAND2X2 U3249 ( .A(n2052), .B(n2053), .Y(n2276) );
  NOR2X4 U3250 ( .A(n2274), .B(n2275), .Y(n2377) );
  NAND2X4 U3251 ( .A(n1897), .B(n3446), .Y(n3445) );
  XOR2X4 U3252 ( .A(n923), .B(n920), .Y(n4078) );
  INVX1 U3253 ( .A(cs[1]), .Y(n2072) );
  INVX4 U3254 ( .A(cs[3]), .Y(n3779) );
  NAND2X4 U3255 ( .A(n571), .B(n577), .Y(n4459) );
  NOR2X2 U3256 ( .A(n1285), .B(n1193), .Y(n1198) );
  NOR2X4 U3257 ( .A(n1141), .B(n1140), .Y(n2055) );
  NAND2X4 U3258 ( .A(n1523), .B(n1524), .Y(n2938) );
  NAND2XL U3259 ( .A(n929), .B(n1094), .Y(n1091) );
  INVXL U3260 ( .A(n929), .Y(n927) );
  OAI22X4 U3261 ( .A0(n1333), .A1(n1956), .B0(n573), .B1(n1955), .Y(n929) );
  AOI21X1 U3262 ( .A0(n3968), .A1(n936), .B0(n3434), .Y(n931) );
  AOI21X4 U3263 ( .A0(n4323), .A1(n968), .B0(n967), .Y(n932) );
  OAI21X4 U3264 ( .A0(n3627), .A1(n958), .B0(n957), .Y(n3898) );
  NOR2X2 U3265 ( .A(n935), .B(n644), .Y(n933) );
  NOR2X4 U3266 ( .A(n1628), .B(n1627), .Y(n4237) );
  INVX2 U3267 ( .A(n3933), .Y(n938) );
  NAND2X2 U3268 ( .A(n1626), .B(n1625), .Y(n3933) );
  INVX4 U3269 ( .A(n1626), .Y(n940) );
  NOR2X4 U3270 ( .A(n4038), .B(n3649), .Y(n943) );
  AOI21X2 U3271 ( .A0(n943), .A1(n3648), .B0(n1872), .Y(n1873) );
  CLKINVX2 U3272 ( .A(n1756), .Y(n945) );
  NAND2X4 U3273 ( .A(n948), .B(n946), .Y(n950) );
  NAND2X4 U3274 ( .A(n950), .B(n1163), .Y(n2849) );
  NAND2X4 U3275 ( .A(n953), .B(n1793), .Y(n1792) );
  NAND2XL U3276 ( .A(n2821), .B(n2822), .Y(n959) );
  OAI21X4 U3277 ( .A0(n3713), .A1(n3712), .B0(n3714), .Y(n1039) );
  NOR2X4 U3278 ( .A(n3415), .B(n3416), .Y(n3713) );
  OR2X4 U3279 ( .A(n2316), .B(n2317), .Y(n2342) );
  INVX2 U3280 ( .A(n2286), .Y(n962) );
  INVX2 U3281 ( .A(n2285), .Y(n963) );
  NAND2BX4 U3282 ( .AN(n2286), .B(n963), .Y(n2337) );
  XNOR2X4 U3283 ( .A(n1223), .B(n1222), .Y(n3237) );
  OAI21X4 U3284 ( .A0(n3594), .A1(n3592), .B0(n3595), .Y(n4323) );
  NOR2X4 U3285 ( .A(n3594), .B(n3591), .Y(n3599) );
  INVXL U3286 ( .A(n970), .Y(n3839) );
  XOR2X1 U3287 ( .A(n971), .B(n973), .Y(n2850) );
  XOR2X1 U3288 ( .A(n972), .B(n974), .Y(n2580) );
  XOR2X1 U3289 ( .A(n971), .B(n975), .Y(n2759) );
  XOR2X2 U3290 ( .A(n972), .B(n590), .Y(n1504) );
  XOR2X1 U3291 ( .A(n971), .B(n1045), .Y(n1600) );
  XOR2X1 U3292 ( .A(n971), .B(n2831), .Y(n2113) );
  XOR2X1 U3293 ( .A(n972), .B(n669), .Y(n1665) );
  XOR2X1 U3294 ( .A(n972), .B(n592), .Y(n2202) );
  XOR2X1 U3295 ( .A(n971), .B(n977), .Y(n2528) );
  XOR2X1 U3296 ( .A(n773), .B(n574), .Y(n2697) );
  XNOR3X2 U3297 ( .A(n2600), .B(n980), .C(n2601), .Y(n2602) );
  OAI22X2 U3298 ( .A0(n2930), .A1(n3091), .B0(n3092), .B1(n986), .Y(n3132) );
  NAND2XL U3299 ( .A(n990), .B(n581), .Y(n989) );
  OAI21X4 U3300 ( .A0(n992), .A1(n4380), .B0(n4381), .Y(n1101) );
  OAI2BB1X2 U3301 ( .A0N(n3038), .A1N(n994), .B0(n993), .Y(n3077) );
  NAND2XL U3302 ( .A(n3039), .B(n996), .Y(n993) );
  NOR2X1 U3303 ( .A(n1337), .B(butt_a_imag[7]), .Y(n1000) );
  NAND2X1 U3304 ( .A(lay_cnt[2]), .B(cs[1]), .Y(n1143) );
  OAI21X4 U3305 ( .A0(n3688), .A1(n3687), .B0(n3689), .Y(n2278) );
  NAND2X2 U3306 ( .A(n1988), .B(n1989), .Y(n3689) );
  NAND2X4 U3307 ( .A(n1987), .B(n1986), .Y(n3687) );
  NOR2X4 U3308 ( .A(n1988), .B(n1989), .Y(n3688) );
  OAI22X2 U3309 ( .A0(n1794), .A1(n2264), .B0(n1755), .B1(n2263), .Y(n1005) );
  OAI22X1 U3310 ( .A0(n2759), .A1(n3068), .B0(n2641), .B1(n3070), .Y(n1009) );
  XOR3X2 U3311 ( .A(n2990), .B(n2989), .C(n2988), .Y(n3001) );
  ADDHX1 U3312 ( .A(n1343), .B(n1342), .CO(n1487), .S(n1346) );
  OAI2BB1X2 U3313 ( .A0N(n2912), .A1N(n3345), .B0(n2911), .Y(n3339) );
  ADDFHX4 U3314 ( .A(n2142), .B(n2141), .CI(n2140), .CO(n2147), .S(n2143) );
  XOR2X1 U3315 ( .A(n593), .B(n1013), .Y(n2752) );
  NAND2X4 U3316 ( .A(n1020), .B(n1019), .Y(n3355) );
  NAND2X2 U3317 ( .A(n3359), .B(n727), .Y(n1019) );
  OAI21X4 U3318 ( .A0(n3359), .A1(n727), .B0(n3358), .Y(n1020) );
  OAI2BB1X4 U3319 ( .A0N(n1023), .A1N(n2988), .B0(n1022), .Y(n3035) );
  NAND2BX2 U3320 ( .AN(n2990), .B(n1024), .Y(n1023) );
  NOR2X4 U3321 ( .A(n2377), .B(n2146), .Y(n2277) );
  NOR2X4 U3322 ( .A(n2052), .B(n2053), .Y(n2146) );
  XOR3X2 U3323 ( .A(n3034), .B(n3035), .C(n3033), .Y(n3063) );
  NAND2X1 U3324 ( .A(n3679), .B(n4537), .Y(n1025) );
  NAND2XL U3325 ( .A(n1469), .B(n1468), .Y(n3679) );
  OAI21X1 U3326 ( .A0(n2017), .A1(n2016), .B0(n2015), .Y(n1029) );
  XOR2X4 U3327 ( .A(n1031), .B(n1271), .Y(n2979) );
  XOR2X1 U3328 ( .A(n2163), .B(n1032), .Y(n2169) );
  XNOR2X4 U3329 ( .A(n1575), .B(n1574), .Y(n2900) );
  NAND2XL U3330 ( .A(n3324), .B(n3323), .Y(n4295) );
  BUFX20 U3331 ( .A(n2937), .Y(n1036) );
  XOR2X1 U3332 ( .A(n1036), .B(n3542), .Y(n3543) );
  XOR2X1 U3333 ( .A(n1036), .B(n3516), .Y(n3517) );
  NAND2X4 U3334 ( .A(n1284), .B(n1077), .Y(n2937) );
  NOR2X4 U3335 ( .A(n2281), .B(n2282), .Y(n4003) );
  XOR2X1 U3336 ( .A(n1038), .B(n1539), .Y(n1377) );
  INVXL U3337 ( .A(n1039), .Y(n3718) );
  AOI21XL U3338 ( .A0(n4376), .A1(n1039), .B0(n4375), .Y(n4377) );
  XOR2X2 U3339 ( .A(n3251), .B(n1041), .Y(n1040) );
  OAI22X1 U3340 ( .A0(n3111), .A1(n3112), .B0(n3110), .B1(n1040), .Y(n3082) );
  NAND2X1 U3341 ( .A(n2824), .B(n2825), .Y(n1042) );
  XNOR3X4 U3342 ( .A(n2825), .B(n1043), .C(n2823), .Y(n2947) );
  INVXL U3343 ( .A(lay_cnt[4]), .Y(n1132) );
  NAND2X4 U3344 ( .A(n2099), .B(lay_cnt[4]), .Y(n1133) );
  OAI22X1 U3345 ( .A0(n3016), .A1(n3177), .B0(n3179), .B1(n1044), .Y(n3062) );
  OAI211X2 U3346 ( .A0(n1281), .A1(n1046), .B0(n1277), .C0(n1278), .Y(n1503)
         );
  INVX4 U3347 ( .A(n1231), .Y(n1046) );
  OAI22X1 U3348 ( .A0(n2568), .A1(n3446), .B0(n3445), .B1(n901), .Y(n1051) );
  XOR2X1 U3349 ( .A(n1038), .B(n572), .Y(n3111) );
  AOI21X4 U3350 ( .A0(n2278), .A1(n2277), .B0(n1055), .Y(n4025) );
  XNOR3X2 U3351 ( .A(n2042), .B(n2044), .C(n2043), .Y(n1057) );
  OAI22X1 U3352 ( .A0(n1106), .A1(n3273), .B0(n3275), .B1(n1058), .Y(n3042) );
  XOR2X1 U3353 ( .A(n3004), .B(n2974), .Y(n3031) );
  XNOR2X4 U3354 ( .A(n1331), .B(butt_b_real[7]), .Y(n2639) );
  XOR3X2 U3355 ( .A(n2869), .B(n2870), .C(n2868), .Y(n2948) );
  NAND2X1 U3356 ( .A(n1067), .B(n844), .Y(n1077) );
  OAI22X2 U3357 ( .A0(n1072), .A1(n3092), .B0(n1070), .B1(n3091), .Y(n2774) );
  NAND2X4 U3358 ( .A(n3414), .B(n3413), .Y(n3712) );
  NAND2X4 U3359 ( .A(n1071), .B(n1231), .Y(n1142) );
  XOR2X1 U3360 ( .A(n2975), .B(n589), .Y(n1072) );
  XOR2X1 U3361 ( .A(n1073), .B(n1045), .Y(n3016) );
  XOR2X2 U3362 ( .A(n1074), .B(n587), .Y(n1559) );
  XOR2X1 U3363 ( .A(n1074), .B(n2005), .Y(n1782) );
  XOR2X1 U3364 ( .A(n1074), .B(n586), .Y(n2180) );
  XOR2X1 U3365 ( .A(n1073), .B(n3516), .Y(n2660) );
  XOR2X2 U3366 ( .A(n1036), .B(n590), .Y(n1084) );
  NAND2X1 U3367 ( .A(n4596), .B(n1086), .Y(n4215) );
  NAND2XL U3368 ( .A(n4594), .B(n1086), .Y(n4204) );
  NAND2XL U3369 ( .A(n4598), .B(n1086), .Y(n4067) );
  OAI22X2 U3370 ( .A0(n3179), .A1(n1652), .B0(n3177), .B1(n1087), .Y(n1719) );
  NOR2X2 U3371 ( .A(n1224), .B(butt_a_imag[4]), .Y(n1089) );
  NAND2X1 U3372 ( .A(n1090), .B(n4594), .Y(n4216) );
  NAND2XL U3373 ( .A(n1090), .B(n4596), .Y(n2333) );
  NAND2XL U3374 ( .A(n1090), .B(n4598), .Y(n4205) );
  NOR2X4 U3375 ( .A(n3413), .B(n3414), .Y(n3721) );
  NAND2XL U3376 ( .A(n2610), .B(n2609), .Y(n1100) );
  NAND2X1 U3377 ( .A(n3420), .B(n3419), .Y(n4381) );
  XOR3X2 U3378 ( .A(n2550), .B(n2548), .C(n2549), .Y(n2607) );
  OAI22X2 U3379 ( .A0(n2977), .A1(n3273), .B0(n3275), .B1(n1106), .Y(n2989) );
  XOR2X2 U3380 ( .A(n2975), .B(n1107), .Y(n1106) );
  ADDFHX1 U3381 ( .A(n2253), .B(n2252), .CI(n2251), .CO(n2296), .S(n2271) );
  ADDFHX1 U3382 ( .A(n1321), .B(n1320), .CI(n1319), .CO(n1502), .S(n1363) );
  ADDFHX4 U3383 ( .A(n1737), .B(n1736), .CI(n1735), .CO(n1742), .S(n1744) );
  ADDFHX4 U3384 ( .A(n1814), .B(n1813), .CI(n1812), .CO(n1818), .S(n1850) );
  XNOR2X1 U3385 ( .A(n3004), .B(n3173), .Y(n1652) );
  ADDFHX4 U3386 ( .A(n1728), .B(n1727), .CI(n1726), .CO(n1733), .S(n1694) );
  AND2X1 U3387 ( .A(n3585), .B(n3584), .Y(n1111) );
  AND2X1 U3388 ( .A(n4005), .B(n4004), .Y(n1114) );
  XOR2XL U3389 ( .A(n3493), .B(n3492), .Y(n1118) );
  AND2X1 U3390 ( .A(n4381), .B(n4382), .Y(n1121) );
  XOR3X2 U3391 ( .A(n1847), .B(n1845), .C(n1846), .Y(n1122) );
  XOR2X1 U3392 ( .A(n4269), .B(n4268), .Y(n1123) );
  XOR2XL U3393 ( .A(n2383), .B(n2069), .Y(n1124) );
  INVXL U3394 ( .A(n1935), .Y(n1932) );
  INVX2 U3395 ( .A(n1217), .Y(n1218) );
  NAND2BXL U3396 ( .AN(n645), .B(n4076), .Y(n2025) );
  XNOR2X1 U3397 ( .A(n579), .B(n4076), .Y(n2530) );
  INVXL U3398 ( .A(n2262), .Y(n2231) );
  INVXL U3399 ( .A(n4085), .Y(n3514) );
  INVXL U3400 ( .A(n3978), .Y(n3485) );
  INVXL U3401 ( .A(n3726), .Y(n3727) );
  INVXL U3402 ( .A(n2084), .Y(n2087) );
  INVXL U3403 ( .A(n3946), .Y(n4247) );
  INVXL U3404 ( .A(n4294), .Y(n4296) );
  XNOR2XL U3405 ( .A(n3981), .B(n3980), .Y(n4525) );
  NOR2X1 U3406 ( .A(n2098), .B(n2090), .Y(n4607) );
  INVXL U3407 ( .A(n4187), .Y(n4569) );
  INVXL U3408 ( .A(n4090), .Y(n4529) );
  XOR2XL U3409 ( .A(n3632), .B(n3631), .Y(n3925) );
  INVXL U3410 ( .A(n4626), .Y(n3853) );
  INVXL U3411 ( .A(n3268), .Y(n3284) );
  INVXL U3412 ( .A(n3266), .Y(n3285) );
  INVXL U3413 ( .A(n1414), .Y(n1424) );
  INVXL U3414 ( .A(n1413), .Y(n1425) );
  NAND2XL U3415 ( .A(Q[1]), .B(n4145), .Y(n1125) );
  INVXL U3416 ( .A(n1126), .Y(n4670) );
  NAND2XL U3417 ( .A(Q[37]), .B(n4145), .Y(n1127) );
  INVXL U3418 ( .A(n1128), .Y(n4672) );
  NAND2XL U3419 ( .A(Q[19]), .B(n4184), .Y(n1129) );
  INVXL U3420 ( .A(n1130), .Y(n4674) );
  NAND2X4 U3421 ( .A(n3752), .B(n3811), .Y(n3851) );
  BUFX2 U3422 ( .A(n1138), .Y(n3840) );
  NOR2X2 U3423 ( .A(n1258), .B(n1135), .Y(n1184) );
  NAND2X4 U3424 ( .A(n1136), .B(n1285), .Y(n1276) );
  NAND3X2 U3425 ( .A(n1143), .B(n1137), .C(n3750), .Y(n1154) );
  NAND4X4 U3426 ( .A(n1153), .B(n1154), .C(n3779), .D(n1139), .Y(n1162) );
  BUFX4 U3427 ( .A(lay_cnt[2]), .Y(n4625) );
  NAND2X1 U3428 ( .A(n1259), .B(n1142), .Y(n1146) );
  NOR2X1 U3429 ( .A(n3750), .B(n3811), .Y(n3789) );
  INVXL U3430 ( .A(n1143), .Y(n1144) );
  NAND4X1 U3431 ( .A(n3789), .B(n1144), .C(lay_cnt[5]), .D(n3779), .Y(n1273)
         );
  INVX2 U3432 ( .A(n1273), .Y(n1215) );
  NAND2X1 U3433 ( .A(n1215), .B(n1276), .Y(n1145) );
  NAND4X2 U3434 ( .A(n1147), .B(n1207), .C(n1146), .D(n1145), .Y(n1148) );
  XOR2X2 U3435 ( .A(n1156), .B(butt_a_imag[6]), .Y(n1158) );
  NOR2X1 U3436 ( .A(n1157), .B(butt_a_imag[5]), .Y(n1149) );
  NAND2X1 U3437 ( .A(n1228), .B(n1220), .Y(n1151) );
  INVX4 U3438 ( .A(n1285), .Y(n1274) );
  XNOR2X1 U3439 ( .A(n3006), .B(n2979), .Y(n1289) );
  XOR2X1 U3440 ( .A(n1157), .B(n1156), .Y(n1159) );
  NOR2X1 U3441 ( .A(n1159), .B(n1158), .Y(n1160) );
  XOR2X1 U3442 ( .A(n1272), .B(n1160), .Y(n1161) );
  NAND2X4 U3443 ( .A(n3106), .B(n1161), .Y(n3109) );
  INVX2 U3444 ( .A(butt_b_imag[3]), .Y(n1225) );
  XNOR2X1 U3445 ( .A(n949), .B(n3253), .Y(n1358) );
  OAI22X1 U3446 ( .A0(n1358), .A1(n3256), .B0(n1237), .B1(n3254), .Y(n1360) );
  NOR2X4 U3447 ( .A(n1276), .B(n1168), .Y(n1169) );
  NOR2BX4 U3448 ( .AN(n1282), .B(n1169), .Y(n1240) );
  INVX2 U3449 ( .A(butt_a_real[4]), .Y(n1179) );
  NAND2X1 U3450 ( .A(n1172), .B(n1171), .Y(n1192) );
  XNOR2X1 U3451 ( .A(n2751), .B(n1192), .Y(n1173) );
  XNOR2X1 U3452 ( .A(n579), .B(n1173), .Y(n1265) );
  INVX2 U3453 ( .A(butt_b_real[4]), .Y(n2744) );
  XOR2X2 U3454 ( .A(n2744), .B(butt_a_real[4]), .Y(n2746) );
  INVX2 U3455 ( .A(butt_a_real[2]), .Y(n1209) );
  NAND2X1 U3456 ( .A(n2897), .B(n1201), .Y(n1177) );
  XOR2X4 U3457 ( .A(n1178), .B(n1177), .Y(n1701) );
  XOR2XL U3458 ( .A(n1182), .B(n2751), .Y(n1183) );
  OAI22XL U3459 ( .A0(n1265), .A1(n1700), .B0(n1322), .B1(n1701), .Y(n1359) );
  INVX2 U3460 ( .A(butt_a_real[7]), .Y(n1331) );
  XNOR2X1 U3461 ( .A(n2639), .B(n1270), .Y(n1190) );
  XOR2XL U3462 ( .A(n1196), .B(n1195), .Y(n1197) );
  NAND2X2 U3463 ( .A(n1198), .B(n1231), .Y(n1354) );
  INVX2 U3464 ( .A(n1234), .Y(n1200) );
  XNOR2X1 U3465 ( .A(n2897), .B(n1201), .Y(n1202) );
  INVX2 U3466 ( .A(butt_a_real[1]), .Y(n1210) );
  XNOR2X2 U3467 ( .A(n1210), .B(butt_b_real[1]), .Y(n2888) );
  NAND2X1 U3468 ( .A(DP_OP_132J1_122_4436_n2999), .B(butt_a_real[0]), .Y(n1242) );
  NAND2X1 U3469 ( .A(n2888), .B(n1242), .Y(n1204) );
  XNOR2X1 U3470 ( .A(n3164), .B(n1606), .Y(n1236) );
  XOR2XL U3471 ( .A(n1210), .B(n1209), .Y(n1211) );
  NAND2X4 U3472 ( .A(n1219), .B(n1218), .Y(n3166) );
  XNOR2X1 U3473 ( .A(n3166), .B(n3173), .Y(n1264) );
  NOR2X1 U3474 ( .A(n1225), .B(butt_a_imag[3]), .Y(n1221) );
  XOR2X1 U3475 ( .A(n1229), .B(n1228), .Y(n1230) );
  NAND2X4 U3476 ( .A(n1235), .B(n1230), .Y(n3177) );
  OAI2BB1X4 U3477 ( .A0N(n1234), .A1N(n1233), .B0(n1232), .Y(n3029) );
  XNOR2X1 U3478 ( .A(n580), .B(n3253), .Y(n1244) );
  BUFX20 U3479 ( .A(n1238), .Y(n3270) );
  OAI22X1 U3480 ( .A0(n1239), .A1(n1793), .B0(n1792), .B1(n587), .Y(n1268) );
  NOR2X4 U3481 ( .A(n1240), .B(n1261), .Y(n2569) );
  XNOR2X1 U3482 ( .A(n3054), .B(n1243), .Y(n1291) );
  XOR2X2 U3483 ( .A(DP_OP_132J1_122_4436_n2999), .B(butt_a_real[0]), .Y(n3275)
         );
  XNOR2X1 U3484 ( .A(n3164), .B(n1243), .Y(n1257) );
  OAI22X1 U3485 ( .A0(n1311), .A1(n3254), .B0(n1244), .B1(n3256), .Y(n1314) );
  XNOR2X1 U3486 ( .A(n725), .B(n1606), .Y(n1312) );
  ADDFX1 U3487 ( .A(n1248), .B(n1247), .CI(n1246), .CO(n1362), .S(n1317) );
  XOR2X2 U3488 ( .A(n1251), .B(butt_a_imag[0]), .Y(n3271) );
  XNOR2X1 U3489 ( .A(n3014), .B(n594), .Y(n1310) );
  NAND2BXL U3490 ( .AN(n645), .B(n3173), .Y(n1254) );
  OAI22X1 U3491 ( .A0(n1254), .A1(n3179), .B0(n3177), .B1(n1045), .Y(n1372) );
  NOR2BX1 U3492 ( .AN(n645), .B(n3179), .Y(n1374) );
  XNOR2X1 U3493 ( .A(n3251), .B(n1173), .Y(n1296) );
  OAI22X1 U3494 ( .A0(n1296), .A1(n1701), .B0(n1255), .B1(n1700), .Y(n1380) );
  XNOR2X1 U3495 ( .A(n3250), .B(n3173), .Y(n1294) );
  OAI22X1 U3496 ( .A0(n1294), .A1(n3179), .B0(n1256), .B1(n3177), .Y(n1379) );
  INVX1 U3497 ( .A(n3818), .Y(n1262) );
  OAI2BB1X4 U3498 ( .A0N(n1262), .A1N(n1261), .B0(n1260), .Y(n3009) );
  XNOR2X1 U3499 ( .A(n3009), .B(n594), .Y(n1279) );
  XNOR2X1 U3500 ( .A(n1038), .B(n1173), .Y(n1297) );
  OAI22XL U3501 ( .A0(n1265), .A1(n1701), .B0(n1297), .B1(n1700), .Y(n1301) );
  ADDFHX1 U3502 ( .A(n1268), .B(n1267), .CI(n1266), .CO(n1352), .S(n1246) );
  NOR2BX2 U3503 ( .AN(n3270), .B(n1956), .Y(n1343) );
  NAND2X1 U3504 ( .A(n1275), .B(n1071), .Y(n1278) );
  OAI2BB1X2 U3505 ( .A0N(n1283), .A1N(n1282), .B0(n1281), .Y(n3010) );
  XNOR2X1 U3506 ( .A(n2976), .B(n1243), .Y(n1290) );
  XNOR2X1 U3507 ( .A(n3270), .B(n1791), .Y(n1286) );
  OAI22X1 U3508 ( .A0(n1793), .A1(n1287), .B0(n1286), .B1(n1792), .Y(n1300) );
  OAI22X1 U3509 ( .A0(n1295), .A1(n3179), .B0(n1294), .B1(n3177), .Y(n1308) );
  ADDFX1 U3510 ( .A(n1303), .B(n1302), .CI(n1301), .CO(n1349), .S(n1304) );
  XNOR2X1 U3511 ( .A(n580), .B(n594), .Y(n1393) );
  XNOR2X1 U3512 ( .A(n3201), .B(n3253), .Y(n1376) );
  OAI22XL U3513 ( .A0(n1312), .A1(n1608), .B0(n1377), .B1(n1607), .Y(n1390) );
  ADDFX1 U3514 ( .A(n1315), .B(n1314), .CI(n1313), .CO(n1318), .S(n1384) );
  OAI22X1 U3515 ( .A0(n1322), .A1(n1700), .B0(n1506), .B1(n1701), .Y(n1512) );
  XNOR2X2 U3516 ( .A(n769), .B(n2979), .Y(n1473) );
  XNOR2X1 U3517 ( .A(n579), .B(n1791), .Y(n1509) );
  XNOR2X1 U3518 ( .A(n3014), .B(n3173), .Y(n1472) );
  INVX2 U3519 ( .A(butt_a_real[8]), .Y(n1330) );
  XNOR2X1 U3520 ( .A(n1482), .B(n2511), .Y(n1329) );
  BUFX4 U3521 ( .A(n1329), .Y(n1954) );
  XOR2X1 U3522 ( .A(n1331), .B(n1330), .Y(n1332) );
  NOR2X2 U3523 ( .A(n645), .B(n572), .Y(n1335) );
  INVX2 U3524 ( .A(n1335), .Y(n1341) );
  XOR2XL U3525 ( .A(n1337), .B(n1336), .Y(n1339) );
  XNOR2X1 U3526 ( .A(n3250), .B(n591), .Y(n1508) );
  XNOR2X1 U3527 ( .A(n3010), .B(n1606), .Y(n1507) );
  OAI22X1 U3528 ( .A0(n1357), .A1(n1607), .B0(n1507), .B1(n1608), .Y(n1493) );
  OAI22X1 U3529 ( .A0(n1358), .A1(n3254), .B0(n1504), .B1(n3256), .Y(n1491) );
  ADDFHX1 U3530 ( .A(n1364), .B(n1363), .CI(n1362), .CO(n1494), .S(n1367) );
  NAND2X2 U3531 ( .A(n3680), .B(n4538), .Y(n1471) );
  ADDHXL U3532 ( .A(n1375), .B(n1374), .CO(n1371), .S(n1440) );
  OAI22XL U3533 ( .A0(n1377), .A1(n1608), .B0(n1408), .B1(n1607), .Y(n1438) );
  ADDFHX1 U3534 ( .A(n1386), .B(n1385), .CI(n1384), .CO(n1369), .S(n1387) );
  ADDFHX1 U3535 ( .A(n1389), .B(n1388), .CI(n1387), .CO(n1463), .S(n1461) );
  ADDFHX1 U3536 ( .A(n1392), .B(n1391), .CI(n1390), .CO(n1385), .S(n1454) );
  BUFX4 U3537 ( .A(n3166), .Y(n3234) );
  OAI22XL U3538 ( .A0(n1412), .A1(n3269), .B0(n1393), .B1(n3271), .Y(n1443) );
  XNOR2X1 U3539 ( .A(n725), .B(n1243), .Y(n1400) );
  OAI22XL U3540 ( .A0(n1400), .A1(n3273), .B0(n1394), .B1(n3275), .Y(n1442) );
  OAI22XL U3541 ( .A0(n1395), .A1(n1608), .B0(n1607), .B1(n1539), .Y(n1403) );
  NAND2BXL U3542 ( .AN(n3239), .B(n3253), .Y(n1396) );
  OAI22XL U3543 ( .A0(n1396), .A1(n3256), .B0(n3254), .B1(n590), .Y(n1402) );
  OAI22XL U3544 ( .A0(n1400), .A1(n3275), .B0(n1406), .B1(n3273), .Y(n1446) );
  ADDHXL U3545 ( .A(n1405), .B(n1404), .CO(n1401), .S(n1422) );
  OAI22XL U3546 ( .A0(n1406), .A1(n3275), .B0(n1415), .B1(n3273), .Y(n1420) );
  OAI22XL U3547 ( .A0(n1408), .A1(n1608), .B0(n1407), .B1(n1607), .Y(n1437) );
  OAI22X1 U3548 ( .A0(n1410), .A1(n3256), .B0(n1409), .B1(n3254), .Y(n1436) );
  OAI22XL U3549 ( .A0(n1412), .A1(n3271), .B0(n1411), .B1(n3269), .Y(n1435) );
  OAI22XL U3550 ( .A0(n1415), .A1(n3275), .B0(n3265), .B1(n3273), .Y(n1423) );
  OAI22XL U3551 ( .A0(n1416), .A1(n3271), .B0(n3239), .B1(n3269), .Y(n1417) );
  ADDFX1 U3552 ( .A(n1422), .B(n1421), .CI(n1420), .CO(n1444), .S(n1427) );
  ADDFX1 U3553 ( .A(n1425), .B(n1424), .CI(n1423), .CO(n1426), .S(n1418) );
  NAND2XL U3554 ( .A(n1431), .B(n1430), .Y(n1432) );
  OAI21X1 U3555 ( .A0(n1434), .A1(n1433), .B0(n1432), .Y(n1451) );
  ADDFHX1 U3556 ( .A(n1440), .B(n1439), .CI(n1438), .CO(n1398), .S(n1456) );
  ADDFX1 U3557 ( .A(n1443), .B(n1442), .CI(n1441), .CO(n1453), .S(n1455) );
  ADDFX1 U3558 ( .A(n1446), .B(n1445), .CI(n1444), .CO(n1447), .S(n1431) );
  AND2X1 U3559 ( .A(n1448), .B(n1447), .Y(n1449) );
  AOI21X1 U3560 ( .A0(n1451), .A1(n1450), .B0(n1449), .Y(n3939) );
  ADDFX1 U3561 ( .A(n1454), .B(n1453), .CI(n1452), .CO(n1460), .S(n1459) );
  NOR2X1 U3562 ( .A(n1459), .B(n1458), .Y(n3936) );
  NAND2XL U3563 ( .A(n1459), .B(n1458), .Y(n3937) );
  OAI21X1 U3564 ( .A0(n3939), .A1(n3936), .B0(n3937), .Y(n4243) );
  NAND2XL U3565 ( .A(n1463), .B(n1462), .Y(n4419) );
  OAI22X1 U3566 ( .A0(n1473), .A1(n3109), .B0(n1544), .B1(n3106), .Y(n1565) );
  NOR2X1 U3567 ( .A(n1519), .B(butt_a_imag[9]), .Y(n1474) );
  NAND2XL U3568 ( .A(n1476), .B(n1475), .Y(n1477) );
  BUFX8 U3569 ( .A(n1524), .Y(n2940) );
  INVXL U3570 ( .A(n1479), .Y(n1480) );
  INVX2 U3571 ( .A(butt_b_real[10]), .Y(n2423) );
  XOR2X2 U3572 ( .A(n2423), .B(butt_a_real[10]), .Y(n2425) );
  NOR2X1 U3573 ( .A(n1530), .B(butt_b_real[9]), .Y(n1481) );
  NAND2X1 U3574 ( .A(n2511), .B(n1482), .Y(n1483) );
  ADDFHX1 U3575 ( .A(n1490), .B(n1489), .CI(n1488), .CO(n1536), .S(n1499) );
  ADDFHX1 U3576 ( .A(n1493), .B(n1492), .CI(n1491), .CO(n1535), .S(n1498) );
  OAI22X1 U3577 ( .A0(n1504), .A1(n3254), .B0(n1525), .B1(n3256), .Y(n1547) );
  OAI22XL U3578 ( .A0(n1516), .A1(n1701), .B0(n1700), .B1(n1506), .Y(n1545) );
  OAI22X1 U3579 ( .A0(n1517), .A1(n3112), .B0(n1508), .B1(n3110), .Y(n1557) );
  OAI22X1 U3580 ( .A0(n1509), .A1(n1792), .B0(n1559), .B1(n1793), .Y(n1556) );
  XOR3X2 U3581 ( .A(n1549), .B(n1548), .C(n1550), .Y(n1570) );
  XOR2XL U3582 ( .A(n1519), .B(n1518), .Y(n1521) );
  NOR2X1 U3583 ( .A(n1521), .B(n1520), .Y(n1522) );
  XOR2X1 U3584 ( .A(n1522), .B(n1575), .Y(n1523) );
  OAI22X2 U3585 ( .A0(n3254), .A1(n1525), .B0(n3256), .B1(n1577), .Y(n1580) );
  INVX2 U3586 ( .A(butt_b_real[11]), .Y(n2437) );
  XNOR2X2 U3587 ( .A(n2437), .B(butt_a_real[11]), .Y(n2435) );
  XNOR2X1 U3588 ( .A(n2435), .B(n1604), .Y(n1528) );
  XOR2X1 U3589 ( .A(n1530), .B(n1529), .Y(n1531) );
  XOR2XL U3590 ( .A(n1532), .B(n2435), .Y(n1533) );
  INVX2 U3591 ( .A(n1528), .Y(n2005) );
  INVXL U3592 ( .A(n1674), .Y(n1579) );
  ADDFHX1 U3593 ( .A(n1537), .B(n1536), .CI(n1535), .CO(n1618), .S(n1567) );
  XNOR2X1 U3594 ( .A(n3270), .B(n1528), .Y(n1541) );
  OAI22X1 U3595 ( .A0(n1543), .A1(n3177), .B0(n1600), .B1(n3179), .Y(n1589) );
  OAI21X1 U3596 ( .A0(n1550), .A1(n1549), .B0(n1548), .Y(n1552) );
  NAND2XL U3597 ( .A(n1550), .B(n1549), .Y(n1551) );
  OAI22X1 U3598 ( .A0(n1559), .A1(n1792), .B0(n1602), .B1(n1793), .Y(n1613) );
  ADDFHX1 U3599 ( .A(n1563), .B(n1562), .CI(n1561), .CO(n1611), .S(n1564) );
  ADDFHX4 U3600 ( .A(n1571), .B(n1572), .CI(n1570), .CO(n1625), .S(n1624) );
  INVX2 U3601 ( .A(butt_b_imag[12]), .Y(n1656) );
  NOR2X1 U3602 ( .A(n1657), .B(butt_a_imag[11]), .Y(n1573) );
  NOR2BX1 U3603 ( .AN(n2569), .B(n2839), .Y(n1676) );
  ADDFHX1 U3604 ( .A(n1581), .B(n1580), .CI(n1579), .CO(n1686), .S(n1594) );
  ADDFHX1 U3605 ( .A(n1584), .B(n1583), .CI(n1582), .CO(n1685), .S(n1587) );
  ADDFHX1 U3606 ( .A(n1590), .B(n1589), .CI(n1588), .CO(n1728), .S(n1586) );
  XNOR2X1 U3607 ( .A(n578), .B(n2979), .Y(n1666) );
  XNOR2X1 U3608 ( .A(n1036), .B(n1173), .Y(n1654) );
  XNOR2X1 U3609 ( .A(n580), .B(n591), .Y(n1672) );
  OAI22X1 U3610 ( .A0(n1593), .A1(n3110), .B0(n1672), .B1(n3112), .Y(n1683) );
  XOR3X2 U3611 ( .A(n1695), .B(n1694), .C(n1696), .Y(n1746) );
  XNOR2X1 U3612 ( .A(n1038), .B(n1528), .Y(n1679) );
  XNOR2X1 U3613 ( .A(n3054), .B(n1791), .Y(n1716) );
  XOR2X2 U3614 ( .A(n2436), .B(butt_a_real[12]), .Y(n2438) );
  NOR2X1 U3615 ( .A(n1634), .B(n681), .Y(n1603) );
  XNOR2X1 U3616 ( .A(n3201), .B(n2900), .Y(n1678) );
  OAI22X1 U3617 ( .A0(n1610), .A1(n1955), .B0(n1677), .B1(n1956), .Y(n1680) );
  ADDFHX4 U3618 ( .A(n1622), .B(n1621), .CI(n1620), .CO(n1627), .S(n1626) );
  XNOR2X1 U3619 ( .A(n2462), .B(n1699), .Y(n1632) );
  XOR2XL U3620 ( .A(n1636), .B(n2462), .Y(n1637) );
  NAND2BX1 U3621 ( .AN(n1719), .B(n1641), .Y(n1645) );
  NAND2X1 U3622 ( .A(n1719), .B(n640), .Y(n1644) );
  OAI2BB1X2 U3623 ( .A0N(n1717), .A1N(n1645), .B0(n1644), .Y(n1811) );
  INVX2 U3624 ( .A(butt_b_imag[14]), .Y(n1766) );
  INVX2 U3625 ( .A(butt_b_imag[13]), .Y(n1767) );
  XNOR2X2 U3626 ( .A(n1767), .B(butt_a_imag[13]), .Y(n1660) );
  NAND2X1 U3627 ( .A(n1660), .B(n1655), .Y(n1649) );
  XOR2X2 U3628 ( .A(n1650), .B(n1649), .Y(n1651) );
  XNOR2X2 U3629 ( .A(n1655), .B(n1660), .Y(n2830) );
  XNOR2X1 U3630 ( .A(n3250), .B(n2830), .Y(n1703) );
  XOR2XL U3631 ( .A(n1657), .B(n1656), .Y(n1659) );
  NOR2X1 U3632 ( .A(n1659), .B(n1658), .Y(n1661) );
  XOR2X1 U3633 ( .A(n1661), .B(n1660), .Y(n1662) );
  NAND2X4 U3634 ( .A(n2839), .B(n1662), .Y(n2836) );
  INVXL U3635 ( .A(n2836), .Y(n1663) );
  OAI2BB2X1 U3636 ( .B0(n1703), .B1(n2839), .A0N(n1664), .A1N(n1663), .Y(n1721) );
  OAI22XL U3637 ( .A0(n3109), .A1(n1666), .B0(n1665), .B1(n3106), .Y(n1720) );
  ADDFHX1 U3638 ( .A(n1669), .B(n1668), .CI(n1667), .CO(n1690), .S(n1731) );
  INVX2 U3639 ( .A(n2830), .Y(n2831) );
  XNOR2X1 U3640 ( .A(n3014), .B(n591), .Y(n1706) );
  OAI22X1 U3641 ( .A0(n1677), .A1(n1955), .B0(n1956), .B1(n1710), .Y(n1709) );
  OAI22XL U3642 ( .A0(n1702), .A1(n2127), .B0(n1679), .B1(n2126), .Y(n1707) );
  ADDFHX1 U3643 ( .A(n1680), .B(n1681), .CI(n1682), .CO(n1693), .S(n1730) );
  ADDFHX1 U3644 ( .A(n1687), .B(n1686), .CI(n1685), .CO(n1691), .S(n1695) );
  ADDFHX4 U3645 ( .A(n1690), .B(n1689), .CI(n1688), .CO(n1816), .S(n1740) );
  NAND2XL U3646 ( .A(n1696), .B(n1695), .Y(n1697) );
  NAND2X1 U3647 ( .A(n1697), .B(n1698), .Y(n1738) );
  XNOR2X1 U3648 ( .A(n3201), .B(n2830), .Y(n1784) );
  OAI22X1 U3649 ( .A0(n1784), .A1(n2839), .B0(n1703), .B1(n2836), .Y(n1808) );
  OAI22XL U3650 ( .A0(n1775), .A1(n3112), .B0(n1706), .B1(n3110), .Y(n1806) );
  XNOR2X1 U3651 ( .A(n2976), .B(n1791), .Y(n1715) );
  OAI22X1 U3652 ( .A0(n1716), .A1(n1792), .B0(n1715), .B1(n1793), .Y(n1725) );
  ADDFHX1 U3653 ( .A(n1722), .B(n1721), .CI(n1720), .CO(n1809), .S(n1723) );
  ADDFHX1 U3654 ( .A(n1731), .B(n1730), .CI(n1729), .CO(n1732), .S(n1737) );
  XOR3X2 U3655 ( .A(n1851), .B(n1850), .C(n1853), .Y(n1861) );
  NOR2X1 U3656 ( .A(n1865), .B(n1864), .Y(n3639) );
  NOR2X2 U3657 ( .A(n3642), .B(n3639), .Y(n3647) );
  XNOR2X2 U3658 ( .A(n1882), .B(butt_b_real[15]), .Y(n2469) );
  XNOR2X1 U3659 ( .A(n2469), .B(n1788), .Y(n1749) );
  XNOR2X1 U3660 ( .A(n3270), .B(n1749), .Y(n1755) );
  OAI21X1 U3661 ( .A0(n1766), .A1(butt_a_imag[14]), .B0(butt_a_imag[13]), .Y(
        n1760) );
  NAND2X1 U3662 ( .A(n1770), .B(n1765), .Y(n1761) );
  INVXL U3663 ( .A(n1762), .Y(n1763) );
  XOR2X1 U3664 ( .A(n1767), .B(n1766), .Y(n1769) );
  NOR2X1 U3665 ( .A(n1769), .B(n1768), .Y(n1771) );
  XOR2X1 U3666 ( .A(n1771), .B(n1770), .Y(n1772) );
  NAND2X4 U3667 ( .A(n2755), .B(n1772), .Y(n2753) );
  OAI22XL U3668 ( .A0(n1775), .A1(n3110), .B0(n1774), .B1(n3112), .Y(n1836) );
  XNOR2X1 U3669 ( .A(n3014), .B(n2900), .Y(n1802) );
  XNOR2X1 U3670 ( .A(n2976), .B(n1954), .Y(n1827) );
  OAI22X1 U3671 ( .A0(n1783), .A1(n1955), .B0(n1827), .B1(n1956), .Y(n1797) );
  OAI22XL U3672 ( .A0(n1829), .A1(n2839), .B0(n1784), .B1(n2836), .Y(n1796) );
  NAND2X1 U3673 ( .A(n1846), .B(n1847), .Y(n1785) );
  INVX2 U3674 ( .A(butt_b_real[16]), .Y(n2451) );
  XOR2X2 U3675 ( .A(n2451), .B(butt_a_real[16]), .Y(n2453) );
  NOR2X1 U3676 ( .A(n1882), .B(butt_b_real[15]), .Y(n1787) );
  NAND2X1 U3677 ( .A(n2469), .B(n1788), .Y(n1789) );
  XNOR2X1 U3678 ( .A(n949), .B(n2900), .Y(n1899) );
  OAI22XL U3679 ( .A0(n1899), .A1(n2940), .B0(n1802), .B1(n2938), .Y(n1915) );
  INVX2 U3680 ( .A(n1822), .Y(n1821) );
  ADDFHX1 U3681 ( .A(n1811), .B(n1810), .CI(n1809), .CO(n1825), .S(n1817) );
  XNOR3X2 U3682 ( .A(n1823), .B(n1821), .C(n1825), .Y(n1857) );
  NAND2X1 U3683 ( .A(n1818), .B(n1857), .Y(n1819) );
  NAND2XL U3684 ( .A(n1822), .B(n1823), .Y(n1824) );
  OAI2BB1X1 U3685 ( .A0N(n1826), .A1N(n1825), .B0(n1824), .Y(n1928) );
  OAI22X1 U3686 ( .A0(n1827), .A1(n1955), .B0(n1890), .B1(n1956), .Y(n1914) );
  XNOR2X1 U3687 ( .A(n3054), .B(n1528), .Y(n1910) );
  OAI22X1 U3688 ( .A0(n1910), .A1(n2127), .B0(n1828), .B1(n2126), .Y(n1913) );
  XNOR2X1 U3689 ( .A(n580), .B(n2830), .Y(n1908) );
  OAI22XL U3690 ( .A0(n1829), .A1(n2836), .B0(n1908), .B1(n2839), .Y(n1912) );
  ADDFHX1 U3691 ( .A(n1834), .B(n1833), .CI(n1832), .CO(n1841), .S(n1810) );
  ADDFHX1 U3692 ( .A(n1838), .B(n1837), .CI(n1836), .CO(n1918), .S(n1839) );
  ADDFHX1 U3693 ( .A(n1841), .B(n1840), .CI(n1839), .CO(n1921), .S(n1849) );
  ADDFHX4 U3694 ( .A(n1844), .B(n1843), .CI(n1842), .CO(n1848), .S(n1851) );
  NAND2X1 U3695 ( .A(n1850), .B(n1851), .Y(n1852) );
  NOR2X4 U3696 ( .A(n1870), .B(n1871), .Y(n4038) );
  OAI21X2 U3697 ( .A0(n3642), .A1(n3640), .B0(n3643), .Y(n3648) );
  NAND2X1 U3698 ( .A(n1869), .B(n1868), .Y(n3650) );
  OAI21X2 U3699 ( .A0(n3650), .A1(n4038), .B0(n4039), .Y(n1872) );
  OAI21X4 U3700 ( .A0(n3638), .A1(n1874), .B0(n1873), .Y(n2349) );
  XNOR2X2 U3701 ( .A(n2409), .B(butt_a_real[17]), .Y(n2455) );
  XOR2X1 U3702 ( .A(n1882), .B(n1881), .Y(n1883) );
  XOR2XL U3703 ( .A(n1884), .B(n2455), .Y(n1885) );
  NAND2X2 U3704 ( .A(n2362), .B(n1885), .Y(n2361) );
  XOR3X2 U3705 ( .A(n1935), .B(n1933), .C(n1936), .Y(n1978) );
  XOR2XL U3706 ( .A(n1893), .B(n1892), .Y(n1895) );
  NOR2X1 U3707 ( .A(n1895), .B(n1894), .Y(n1896) );
  XOR2XL U3708 ( .A(n1896), .B(n1940), .Y(n1897) );
  XNOR2X1 U3709 ( .A(n579), .B(n1749), .Y(n1958) );
  NAND2BX1 U3710 ( .AN(n3270), .B(n1880), .Y(n1906) );
  OAI22X2 U3711 ( .A0(n1906), .A1(n2362), .B0(n2361), .B1(n586), .Y(n1960) );
  XNOR2X1 U3712 ( .A(n3014), .B(n2830), .Y(n1961) );
  OAI22X1 U3713 ( .A0(n1908), .A1(n2836), .B0(n1961), .B1(n2839), .Y(n1974) );
  XNOR2X1 U3714 ( .A(n2976), .B(n1528), .Y(n1971) );
  OAI22X1 U3715 ( .A0(n1910), .A1(n2126), .B0(n1971), .B1(n2127), .Y(n1963) );
  INVX2 U3716 ( .A(butt_a_imag[18]), .Y(n3530) );
  NOR2BX1 U3717 ( .AN(n645), .B(n4078), .Y(n1994) );
  INVXL U3718 ( .A(n1941), .Y(n1942) );
  ADDFHX1 U3719 ( .A(n1945), .B(n1946), .CI(n1944), .CO(n2043), .S(n1977) );
  INVX2 U3720 ( .A(butt_b_real[18]), .Y(n1998) );
  XOR2X1 U3721 ( .A(n3488), .B(n1998), .Y(n2411) );
  XNOR2X1 U3722 ( .A(n2411), .B(n1950), .Y(n1953) );
  NAND2X1 U3723 ( .A(n2455), .B(n1951), .Y(n1952) );
  XOR2X4 U3724 ( .A(n1953), .B(n1952), .Y(n3558) );
  OAI22XL U3725 ( .A0(n1958), .A1(n2263), .B0(n2027), .B1(n2264), .Y(n2019) );
  ADDFX1 U3726 ( .A(n1964), .B(n1963), .CI(n1962), .CO(n2015), .S(n1947) );
  ADDFHX4 U3727 ( .A(n1967), .B(n1966), .CI(n1965), .CO(n2050), .S(n1984) );
  ADDFHX1 U3728 ( .A(n1970), .B(n1969), .CI(n1968), .CO(n2032), .S(n1967) );
  XNOR2X1 U3729 ( .A(n1036), .B(n1528), .Y(n2006) );
  OAI22X1 U3730 ( .A0(n1971), .A1(n2126), .B0(n2006), .B1(n2127), .Y(n2038) );
  XNOR2X1 U3731 ( .A(n3054), .B(n2197), .Y(n2028) );
  OAI22X1 U3732 ( .A0(n2028), .A1(n2199), .B0(n1972), .B1(n2198), .Y(n2037) );
  ADDFHX4 U3733 ( .A(n1974), .B(n1975), .CI(n1976), .CO(n2034), .S(n1948) );
  ADDFHX4 U3734 ( .A(n1985), .B(n1984), .CI(n1983), .CO(n1989), .S(n1987) );
  INVXL U3735 ( .A(n2372), .Y(n1991) );
  INVXL U3736 ( .A(n2278), .Y(n1990) );
  ADDFHX1 U3737 ( .A(n1994), .B(n1993), .CI(n1992), .CO(n2134), .S(n2044) );
  NAND2X4 U3738 ( .A(n3558), .B(n2003), .Y(n3557) );
  NAND2X1 U3739 ( .A(n2008), .B(n2007), .Y(n3516) );
  XNOR2X1 U3740 ( .A(n3250), .B(n4076), .Y(n2116) );
  XOR2XL U3741 ( .A(butt_b_imag[18]), .B(n2009), .Y(n2011) );
  NAND2X4 U3742 ( .A(n4078), .B(n2012), .Y(n4077) );
  OAI22XL U3743 ( .A0(n2116), .A1(n4078), .B0(n2013), .B1(n4077), .Y(n2111) );
  OAI22XL U3744 ( .A0(n2014), .A1(n2836), .B0(n2113), .B1(n2839), .Y(n2110) );
  NAND2XL U3745 ( .A(n2017), .B(n2016), .Y(n2018) );
  ADDFHX1 U3746 ( .A(n2021), .B(n2020), .CI(n2019), .CO(n2124), .S(n2016) );
  XNOR2X1 U3747 ( .A(n579), .B(n1880), .Y(n2128) );
  XNOR2X1 U3748 ( .A(n2976), .B(n2197), .Y(n2125) );
  XNOR2X1 U3749 ( .A(n769), .B(n2567), .Y(n2118) );
  ADDFHX4 U3750 ( .A(n2031), .B(n2032), .CI(n2030), .CO(n2144), .S(n2049) );
  ADDFHX1 U3751 ( .A(n2041), .B(n2040), .CI(n2039), .CO(n2136), .S(n2017) );
  NAND2XL U3752 ( .A(n2042), .B(n2044), .Y(n2046) );
  OAI21X1 U3753 ( .A0(n2042), .A1(n2044), .B0(n2043), .Y(n2045) );
  NAND2X1 U3754 ( .A(n2046), .B(n2045), .Y(n2135) );
  NAND2X1 U3755 ( .A(Q[0]), .B(butt_a_imag[0]), .Y(n3944) );
  OAI21X1 U3756 ( .A0(n3941), .A1(n3944), .B0(n3942), .Y(n3946) );
  OAI21XL U3757 ( .A0(n4248), .A1(n4245), .B0(n4249), .Y(n2058) );
  NAND2XL U3758 ( .A(n3658), .B(n2061), .Y(n2063) );
  OAI21XL U3759 ( .A0(n3668), .A1(n3664), .B0(n3669), .Y(n3657) );
  NAND2XL U3760 ( .A(Q[6]), .B(butt_a_imag[6]), .Y(n4051) );
  OAI21XL U3761 ( .A0(n4054), .A1(n4051), .B0(n4055), .Y(n2060) );
  AOI21XL U3762 ( .A0(n2061), .A1(n3657), .B0(n2060), .Y(n2062) );
  NAND2XL U3763 ( .A(n2084), .B(n2065), .Y(n4044) );
  OAI21XL U3764 ( .A0(n3695), .A1(n3701), .B0(n3696), .Y(n2085) );
  OAI21XL U3765 ( .A0(n2389), .A1(n2385), .B0(n2390), .Y(n2064) );
  AOI21XL U3766 ( .A0(n2065), .A1(n2085), .B0(n2064), .Y(n4043) );
  OAI21XL U3767 ( .A0(n4043), .A1(n4046), .B0(n4047), .Y(n2066) );
  INVXL U3768 ( .A(n2074), .Y(n2068) );
  AOI21X1 U3769 ( .A0(n2077), .A1(n2075), .B0(n2068), .Y(n2097) );
  NAND2XL U3770 ( .A(Q[15]), .B(butt_a_imag[15]), .Y(n2094) );
  OAI21X1 U3771 ( .A0(n2097), .A1(n2093), .B0(n2094), .Y(n2383) );
  NAND2XL U3772 ( .A(n2382), .B(n2380), .Y(n2069) );
  NAND2X2 U3773 ( .A(n4111), .B(n4184), .Y(n2098) );
  NOR2X1 U3774 ( .A(n2098), .B(n4502), .Y(n2071) );
  NAND2XL U3775 ( .A(n2075), .B(n2074), .Y(n2076) );
  NOR4XL U3776 ( .A(in_out_cnt[4]), .B(in_out_cnt[3]), .C(in_out_cnt[2]), .D(
        in_out_cnt[0]), .Y(n2078) );
  INVXL U3777 ( .A(in_out_cnt[10]), .Y(n4665) );
  INVXL U3778 ( .A(in_out_cnt[1]), .Y(n4631) );
  NAND4XL U3779 ( .A(n2078), .B(n4665), .C(n4647), .D(n4631), .Y(n2080) );
  INVXL U3780 ( .A(in_out_cnt[8]), .Y(n4636) );
  INVXL U3781 ( .A(in_out_cnt[6]), .Y(n3845) );
  NAND4XL U3782 ( .A(n4636), .B(n3833), .C(n3845), .D(n3837), .Y(n2079) );
  INVXL U3783 ( .A(n2085), .Y(n2086) );
  INVXL U3784 ( .A(n2088), .Y(n2387) );
  NAND2XL U3785 ( .A(n2387), .B(n2385), .Y(n2089) );
  AOI22XL U3786 ( .A0(n4608), .A1(FFT2D_IN_R[14]), .B0(n4604), .B1(n4607), .Y(
        n2091) );
  OAI2BB1XL U3787 ( .A0N(FFT2D_IN_I[14]), .A1N(n4600), .B0(n2091), .Y(n2092)
         );
  AOI21XL U3788 ( .A0(n4602), .A1(n4208), .B0(n2092), .Y(n2104) );
  INVXL U3789 ( .A(n2093), .Y(n2095) );
  NAND2XL U3790 ( .A(n2095), .B(n2094), .Y(n2096) );
  XOR2X1 U3791 ( .A(n2097), .B(n2096), .Y(n4206) );
  INVXL U3792 ( .A(n4234), .Y(n2102) );
  NAND2XL U3793 ( .A(n4206), .B(n4605), .Y(n2103) );
  OAI211X1 U3794 ( .A0(n1124), .A1(n4552), .B0(n2104), .C0(n2103), .Y(n2105)
         );
  ADDHX1 U3795 ( .A(n2106), .B(n2107), .CO(n2160), .S(n2130) );
  ADDFHX1 U3796 ( .A(n2111), .B(n2112), .CI(n2110), .CO(n2158), .S(n2132) );
  OAI22X1 U3797 ( .A0(n2113), .A1(n2836), .B0(n2161), .B1(n2839), .Y(n2167) );
  XNOR2X1 U3798 ( .A(n3201), .B(n4076), .Y(n2179) );
  OAI22XL U3799 ( .A0(n2118), .A1(n3445), .B0(n2182), .B1(n3446), .Y(n2174) );
  ADDFHX1 U3800 ( .A(n2121), .B(n2120), .CI(n2119), .CO(n2171), .S(n2122) );
  OAI22XL U3801 ( .A0(n2128), .A1(n2361), .B0(n2180), .B1(n2362), .Y(n2168) );
  ADDFHX1 U3802 ( .A(n2129), .B(n2130), .CI(n2131), .CO(n2184), .S(n2123) );
  ADDFHX4 U3803 ( .A(n2149), .B(n2147), .CI(n2148), .CO(n2279), .S(n2274) );
  OAI2BB1X2 U3804 ( .A0N(n2157), .A1N(n2156), .B0(n2155), .Y(n2188) );
  ADDFX1 U3805 ( .A(n2160), .B(n2159), .CI(n2158), .CO(n2192), .S(n2152) );
  XNOR2X1 U3806 ( .A(n3004), .B(n2830), .Y(n2200) );
  ADDFHX1 U3807 ( .A(n2166), .B(n2167), .CI(n2165), .CO(n2220), .S(n2173) );
  ADDFHX1 U3808 ( .A(n2173), .B(n2171), .CI(n2172), .CO(n2190), .S(n2151) );
  ADDFHX1 U3809 ( .A(n2176), .B(n2175), .CI(n2174), .CO(n2210), .S(n2172) );
  XNOR2X1 U3810 ( .A(n579), .B(n3556), .Y(n2205) );
  XNOR2X1 U3811 ( .A(n769), .B(n4076), .Y(n2215) );
  OAI22XL U3812 ( .A0(n2215), .A1(n4078), .B0(n2179), .B1(n4077), .Y(n2206) );
  OAI22XL U3813 ( .A0(n2180), .A1(n2361), .B0(n2362), .B1(n2204), .Y(n2213) );
  OAI22X1 U3814 ( .A0(n2181), .A1(n2263), .B0(n2203), .B1(n2264), .Y(n2212) );
  BUFX2 U3815 ( .A(n3014), .Y(n2675) );
  XNOR2X1 U3816 ( .A(n2675), .B(n2567), .Y(n2214) );
  OAI22XL U3817 ( .A0(n2182), .A1(n3445), .B0(n2214), .B1(n3446), .Y(n2211) );
  ADDFHX4 U3818 ( .A(n2185), .B(n2184), .CI(n2183), .CO(n2194), .S(n2153) );
  INVXL U3819 ( .A(n2200), .Y(n2201) );
  OAI2BB1X1 U3820 ( .A0N(n2839), .A1N(n2836), .B0(n2201), .Y(n2230) );
  OAI22X1 U3821 ( .A0(n2203), .A1(n2263), .B0(n2233), .B1(n2264), .Y(n2239) );
  OAI22XL U3822 ( .A0(n2205), .A1(n3557), .B0(n2228), .B1(n3558), .Y(n2237) );
  ADDFX1 U3823 ( .A(n2213), .B(n2212), .CI(n2211), .CO(n2227), .S(n2208) );
  BUFX2 U3824 ( .A(n949), .Y(n2700) );
  XNOR2X1 U3825 ( .A(n2700), .B(n2567), .Y(n2242) );
  OAI22XL U3826 ( .A0(n2215), .A1(n4077), .B0(n2240), .B1(n4078), .Y(n2244) );
  ADDFHX1 U3827 ( .A(n2218), .B(n2217), .CI(n2216), .CO(n2243), .S(n2221) );
  OAI22XL U3828 ( .A0(n2228), .A1(n3557), .B0(n2269), .B1(n3558), .Y(n2259) );
  ADDFHX1 U3829 ( .A(n2231), .B(n2230), .CI(n2229), .CO(n2258), .S(n2236) );
  ADDFX1 U3830 ( .A(n2245), .B(n2244), .CI(n2243), .CO(n2251), .S(n2226) );
  ADDFHX1 U3831 ( .A(n2259), .B(n2258), .CI(n2257), .CO(n2312), .S(n2273) );
  OAI2BB1X1 U3832 ( .A0N(n2264), .A1N(n2263), .B0(n1749), .Y(n2359) );
  OAI2BB1X1 U3833 ( .A0N(n2755), .A1N(n2753), .B0(n2266), .Y(n2308) );
  XNOR2X1 U3834 ( .A(n1036), .B(n1880), .Y(n2301) );
  XNOR2X1 U3835 ( .A(n3054), .B(n3556), .Y(n2306) );
  OAI22X1 U3836 ( .A0(n2306), .A1(n3558), .B0(n2269), .B1(n3557), .Y(n2303) );
  XNOR2X1 U3837 ( .A(n2700), .B(n4076), .Y(n2305) );
  XNOR3X2 U3838 ( .A(n2310), .B(n2312), .C(n2314), .Y(n2295) );
  NAND2X1 U3839 ( .A(n595), .B(n2337), .Y(n2289) );
  INVX3 U3840 ( .A(n4025), .Y(n4000) );
  INVX1 U3841 ( .A(n2346), .Y(n2320) );
  NAND2X1 U3842 ( .A(n2284), .B(n2283), .Y(n2344) );
  INVXL U3843 ( .A(n2344), .Y(n2287) );
  AOI21XL U3844 ( .A0(n2287), .A1(n2337), .B0(n2343), .Y(n2288) );
  AOI21X1 U3845 ( .A0(n4000), .A1(n2291), .B0(n2290), .Y(n2292) );
  ADDFHX1 U3846 ( .A(n2299), .B(n2298), .CI(n2297), .CO(n2352), .S(n2314) );
  ADDFX1 U3847 ( .A(n2304), .B(n2303), .CI(n2302), .CO(n2367), .S(n2297) );
  XNOR2X1 U3848 ( .A(n773), .B(n4076), .Y(n2365) );
  XNOR2X1 U3849 ( .A(n2976), .B(n3556), .Y(n2356) );
  NAND2XL U3850 ( .A(n2312), .B(n2311), .Y(n2313) );
  NAND2XL U3851 ( .A(n2317), .B(n2316), .Y(n2340) );
  NAND2X1 U3852 ( .A(n2342), .B(n2340), .Y(n2318) );
  NAND2XL U3853 ( .A(n4230), .B(n4598), .Y(n2335) );
  OAI21X1 U3854 ( .A0(n2320), .A1(n2338), .B0(n2344), .Y(n2321) );
  AOI21X1 U3855 ( .A0(n4000), .A1(n2322), .B0(n2321), .Y(n2323) );
  OAI21X2 U3856 ( .A0(n2324), .A1(n4027), .B0(n2323), .Y(n2327) );
  NAND2X1 U3857 ( .A(n2325), .B(n2337), .Y(n2326) );
  NOR2X4 U3858 ( .A(n2371), .B(n4234), .Y(n4594) );
  NAND2X1 U3859 ( .A(n3998), .B(n2339), .Y(n2329) );
  ADDFX1 U3860 ( .A(n2355), .B(n2354), .CI(n2353), .CO(n3537), .S(n2366) );
  ADDFX1 U3861 ( .A(n2359), .B(n2358), .CI(n2357), .CO(n3545), .S(n2368) );
  INVXL U3862 ( .A(n2363), .Y(n2364) );
  ADDFX1 U3863 ( .A(n2368), .B(n2367), .CI(n2366), .CO(n3535), .S(n2351) );
  INVXL U3864 ( .A(n2276), .Y(n2373) );
  INVXL U3865 ( .A(n2380), .Y(n2381) );
  INVXL U3866 ( .A(n2385), .Y(n2386) );
  INVXL U3867 ( .A(n2389), .Y(n2391) );
  NAND2XL U3868 ( .A(n2391), .B(n2390), .Y(n2392) );
  AOI22XL U3869 ( .A0(n4600), .A1(FFT2D_IN_I[15]), .B0(FFT2D_IN_R[15]), .B1(
        n4608), .Y(n2394) );
  OAI2BB1XL U3870 ( .A0N(n4607), .A1N(n4601), .B0(n2394), .Y(n2395) );
  XNOR2X1 U3871 ( .A(n2411), .B(n2404), .Y(n2408) );
  NAND2X1 U3872 ( .A(n2455), .B(n2445), .Y(n2407) );
  XOR2XL U3873 ( .A(butt_b_real[18]), .B(n2409), .Y(n2410) );
  NAND2X2 U3874 ( .A(n4082), .B(n2412), .Y(n4081) );
  OAI22X1 U3875 ( .A0(n2414), .A1(n4082), .B0(n4081), .B1(n2413), .Y(n2495) );
  OAI21X1 U3876 ( .A0(n2423), .A1(butt_a_real[10]), .B0(butt_a_real[9]), .Y(
        n2417) );
  NAND2XL U3877 ( .A(butt_a_real[10]), .B(n2423), .Y(n2416) );
  NAND2X1 U3878 ( .A(n2417), .B(n2416), .Y(n2434) );
  NOR2X1 U3879 ( .A(n2424), .B(butt_a_real[9]), .Y(n2418) );
  NAND2X1 U3880 ( .A(n2511), .B(n2510), .Y(n2421) );
  XOR2XL U3881 ( .A(n2424), .B(n2423), .Y(n2426) );
  NOR2X1 U3882 ( .A(n2426), .B(n2425), .Y(n2427) );
  XOR2XL U3883 ( .A(n2427), .B(n2435), .Y(n2428) );
  NAND2X2 U3884 ( .A(n3087), .B(n2428), .Y(n3085) );
  XOR2XL U3885 ( .A(n2440), .B(n2462), .Y(n2441) );
  NAND2X2 U3886 ( .A(n2883), .B(n2441), .Y(n2846) );
  OAI22XL U3887 ( .A0(n2571), .A1(n2846), .B0(n2883), .B1(n2442), .Y(n2518) );
  OAI22X1 U3888 ( .A0(n2490), .A1(n2755), .B0(n2444), .B1(n2753), .Y(n2476) );
  XNOR2X1 U3889 ( .A(n2976), .B(n2830), .Y(n2480) );
  OAI22X1 U3890 ( .A0(n2564), .A1(n2836), .B0(n2480), .B1(n2839), .Y(n2558) );
  XNOR2X2 U3891 ( .A(n2455), .B(n2445), .Y(n2711) );
  NOR2X1 U3892 ( .A(n2452), .B(butt_a_real[15]), .Y(n2446) );
  NAND2X1 U3893 ( .A(n2448), .B(n2447), .Y(n2459) );
  XOR2XL U3894 ( .A(n2452), .B(n2451), .Y(n2454) );
  NOR2X1 U3895 ( .A(n2454), .B(n733), .Y(n2456) );
  XOR2XL U3896 ( .A(n2456), .B(n2455), .Y(n2457) );
  NAND2X2 U3897 ( .A(n3450), .B(n2457), .Y(n3449) );
  NOR2X1 U3898 ( .A(n2466), .B(butt_a_real[13]), .Y(n2460) );
  NAND2X1 U3899 ( .A(n2462), .B(n2461), .Y(n2463) );
  XOR2X1 U3900 ( .A(n2466), .B(n2465), .Y(n2468) );
  NOR2X1 U3901 ( .A(n2468), .B(n2467), .Y(n2470) );
  XOR2XL U3902 ( .A(n2470), .B(n2469), .Y(n2471) );
  NAND2X4 U3903 ( .A(n2765), .B(n2471), .Y(n2763) );
  OAI22X1 U3904 ( .A0(n2486), .A1(n2765), .B0(n2497), .B1(n2763), .Y(n2484) );
  OAI22XL U3905 ( .A0(n2479), .A1(n2836), .B0(n2839), .B1(n2831), .Y(n2541) );
  OAI22XL U3906 ( .A0(n2836), .A1(n2480), .B0(n2479), .B1(n2839), .Y(n2494) );
  XNOR2X1 U3907 ( .A(n2481), .B(n2482), .Y(n2493) );
  OAI22XL U3908 ( .A0(n2498), .A1(n3445), .B0(n2489), .B1(n3446), .Y(n2492) );
  ADDFHX1 U3909 ( .A(n2485), .B(n2484), .CI(n2483), .CO(n2535), .S(n2551) );
  OAI22X1 U3910 ( .A0(n2540), .A1(n4082), .B0(n4081), .B1(n2488), .Y(n2531) );
  OAI22X1 U3911 ( .A0(n2490), .A1(n2753), .B0(n2529), .B1(n2755), .Y(n2537) );
  ADDFHX1 U3912 ( .A(n2494), .B(n2493), .CI(n2492), .CO(n2544), .S(n2583) );
  ADDHX1 U3913 ( .A(n2496), .B(n2495), .CO(n2550), .S(n2562) );
  OAI22X1 U3914 ( .A0(n2565), .A1(n2763), .B0(n2497), .B1(n2765), .Y(n2561) );
  XOR2X4 U3915 ( .A(n2503), .B(n2502), .Y(n3070) );
  XOR2XL U3916 ( .A(n2505), .B(n2504), .Y(n2507) );
  NOR2X1 U3917 ( .A(n2507), .B(n2506), .Y(n2508) );
  XOR2XL U3918 ( .A(n2508), .B(n2511), .Y(n2509) );
  XNOR2X1 U3919 ( .A(n2511), .B(n2510), .Y(n2512) );
  INVXL U3920 ( .A(n2572), .Y(n2513) );
  OAI2BB1X1 U3921 ( .A0N(n3070), .A1N(n3068), .B0(n2513), .Y(n2576) );
  OAI2BB1X4 U3922 ( .A0N(n2601), .A1N(n2525), .B0(n2524), .Y(n2726) );
  OAI2BB1X1 U3923 ( .A0N(n2883), .A1N(n2846), .B0(n2527), .Y(n2662) );
  XNOR2X1 U3924 ( .A(n1036), .B(n657), .Y(n2665) );
  XNOR2X1 U3925 ( .A(n3054), .B(n2567), .Y(n2673) );
  OAI22X1 U3926 ( .A0(n2530), .A1(n4077), .B0(n2660), .B1(n4078), .Y(n2669) );
  ADDFHX1 U3927 ( .A(n2535), .B(n2533), .CI(n2534), .CO(n2681), .S(n2599) );
  INVX1 U3928 ( .A(n2655), .Y(n2547) );
  XNOR2X1 U3929 ( .A(n949), .B(n2711), .Y(n2672) );
  OAI22X1 U3930 ( .A0(n2540), .A1(n4081), .B0(n2676), .B1(n4082), .Y(n2678) );
  ADDFHX1 U3931 ( .A(n2543), .B(n2542), .CI(n2541), .CO(n2677), .S(n2546) );
  XNOR3X2 U3932 ( .A(n2547), .B(n2656), .C(n2658), .Y(n2680) );
  OAI22X1 U3933 ( .A0(n2618), .A1(n2753), .B0(n2755), .B1(n2556), .Y(n2587) );
  XNOR2X1 U3934 ( .A(n2976), .B(n2900), .Y(n2594) );
  OAI22X1 U3935 ( .A0(n2594), .A1(n2938), .B0(n2563), .B1(n2940), .Y(n2625) );
  XNOR2X1 U3936 ( .A(n3164), .B(n2830), .Y(n2593) );
  OAI22X1 U3937 ( .A0(n2564), .A1(n2839), .B0(n2593), .B1(n2836), .Y(n2624) );
  XNOR2X1 U3938 ( .A(n3234), .B(n2757), .Y(n2595) );
  OAI22X1 U3939 ( .A0(n2566), .A1(n3450), .B0(n2579), .B1(n3449), .Y(n2592) );
  NAND2BXL U3940 ( .AN(n2569), .B(n2711), .Y(n2570) );
  OAI22XL U3941 ( .A0(n2571), .A1(n2883), .B0(n2617), .B1(n2846), .Y(n2590) );
  XNOR2X1 U3942 ( .A(n2975), .B(n2512), .Y(n2641) );
  OAI22X1 U3943 ( .A0(n2641), .A1(n3068), .B0(n2572), .B1(n3070), .Y(n2643) );
  XNOR2X1 U3944 ( .A(n3265), .B(n2567), .Y(n2573) );
  OAI22X1 U3945 ( .A0(n2574), .A1(n3446), .B0(n2573), .B1(n3445), .Y(n2642) );
  OAI22X1 U3946 ( .A0(n2579), .A1(n3450), .B0(n2578), .B1(n3449), .Y(n2646) );
  XNOR2X1 U3947 ( .A(n949), .B(n3084), .Y(n2770) );
  ADDFHX1 U3948 ( .A(n2592), .B(n2591), .CI(n2590), .CO(n2649), .S(n2612) );
  OAI22XL U3949 ( .A0(n2616), .A1(n2836), .B0(n2593), .B1(n2839), .Y(n2622) );
  XNOR2X1 U3950 ( .A(n3054), .B(n2900), .Y(n2734) );
  OAI22X1 U3951 ( .A0(n2734), .A1(n2938), .B0(n2594), .B1(n2940), .Y(n2621) );
  ADDFHX4 U3952 ( .A(n2613), .B(n639), .CI(n2611), .CO(n2954), .S(n2732) );
  XNOR2X1 U3953 ( .A(n2615), .B(n2614), .Y(n2804) );
  XNOR2X1 U3954 ( .A(n579), .B(n2830), .Y(n2738) );
  XNOR2X1 U3955 ( .A(n3029), .B(n2432), .Y(n2735) );
  NOR2BX1 U3956 ( .AN(n3239), .B(n3450), .Y(n2772) );
  NOR2X1 U3957 ( .A(n2635), .B(butt_a_real[5]), .Y(n2631) );
  OAI21X1 U3958 ( .A0(butt_a_real[4]), .A1(n2744), .B0(butt_a_real[3]), .Y(
        n2633) );
  XOR2X1 U3959 ( .A(n2635), .B(n2634), .Y(n2636) );
  XOR2XL U3960 ( .A(n2637), .B(n2639), .Y(n2638) );
  NAND2X2 U3961 ( .A(n3091), .B(n2638), .Y(n3092) );
  ADDFHX1 U3962 ( .A(n2647), .B(n2646), .CI(n2645), .CO(n2608), .S(n2811) );
  ADDFHX4 U3963 ( .A(n2654), .B(n2653), .CI(n2652), .CO(n2603), .S(n2962) );
  NAND2XL U3964 ( .A(n2656), .B(n2655), .Y(n2657) );
  OAI2BB1X1 U3965 ( .A0N(n2658), .A1N(n2659), .B0(n2657), .Y(n2730) );
  XNOR2X1 U3966 ( .A(n3164), .B(n4076), .Y(n2699) );
  ADDFHX1 U3967 ( .A(n2663), .B(n2662), .CI(n2661), .CO(n2690), .S(n2668) );
  ADDFX1 U3968 ( .A(n2669), .B(n2670), .CI(n2671), .CO(n2685), .S(n2667) );
  OAI22X1 U3969 ( .A0(n2672), .A1(n3449), .B0(n2697), .B1(n3450), .Y(n2688) );
  XNOR2X1 U3970 ( .A(n2675), .B(n2674), .Y(n2701) );
  OAI22XL U3971 ( .A0(n2676), .A1(n4081), .B0(n2701), .B1(n4082), .Y(n2686) );
  ADDFHX1 U3972 ( .A(n2685), .B(n2684), .CI(n2683), .CO(n2707), .S(n2702) );
  XNOR2X1 U3973 ( .A(n1036), .B(n2567), .Y(n2713) );
  XNOR2X1 U3974 ( .A(n3054), .B(n4076), .Y(n2718) );
  XNOR2X1 U3975 ( .A(n2700), .B(n2674), .Y(n2717) );
  ADDFHX4 U3976 ( .A(n2704), .B(n2703), .CI(n2702), .CO(n2705), .S(n2729) );
  ADDFX1 U3977 ( .A(n2716), .B(n2715), .CI(n2714), .CO(n3454), .S(n2708) );
  XNOR2X1 U3978 ( .A(n773), .B(n2674), .Y(n3452) );
  XNOR2X1 U3979 ( .A(n2733), .B(n2900), .Y(n2790) );
  XNOR2X1 U3980 ( .A(n3014), .B(n3084), .Y(n2769) );
  XNOR2X1 U3981 ( .A(n3029), .B(n3084), .Y(n2828) );
  NOR2BX1 U3982 ( .AN(n645), .B(n2765), .Y(n2844) );
  NOR2X1 U3983 ( .A(n2745), .B(butt_a_real[3]), .Y(n2739) );
  INVX2 U3984 ( .A(butt_b_real[2]), .Y(n2891) );
  NAND2X1 U3985 ( .A(n2897), .B(n2896), .Y(n2742) );
  XOR2XL U3986 ( .A(n2745), .B(n2744), .Y(n2747) );
  NOR2X1 U3987 ( .A(n2747), .B(n2746), .Y(n2748) );
  XOR2XL U3988 ( .A(n2748), .B(n2751), .Y(n2749) );
  NAND2X2 U3989 ( .A(n3184), .B(n2749), .Y(n3182) );
  OAI22X1 U3990 ( .A0(n2834), .A1(n3068), .B0(n2759), .B1(n3070), .Y(n2776) );
  ADDFHX1 U3991 ( .A(n2762), .B(n2761), .CI(n2760), .CO(n2808), .S(n2825) );
  NAND2XL U3992 ( .A(n2794), .B(n2795), .Y(n2779) );
  NAND2X1 U3993 ( .A(n2780), .B(n2779), .Y(n2806) );
  XNOR2X1 U3994 ( .A(n2782), .B(n2781), .Y(n2859) );
  XNOR2X1 U3995 ( .A(n2783), .B(n2830), .Y(n2838) );
  XNOR2X1 U3996 ( .A(n579), .B(n2900), .Y(n2860) );
  OAI22X1 U3997 ( .A0(n2860), .A1(n2938), .B0(n2791), .B1(n2940), .Y(n2857) );
  ADDFHX1 U3998 ( .A(n2801), .B(n2799), .CI(n2800), .CO(n2807), .S(n2815) );
  ADDFHX4 U3999 ( .A(n2816), .B(n2815), .CI(n2814), .CO(n2821), .S(n2872) );
  XNOR2X1 U4000 ( .A(n2976), .B(n2979), .Y(n2905) );
  XNOR2X1 U4001 ( .A(n769), .B(n3084), .Y(n2861) );
  OAI22XL U4002 ( .A0(n2861), .A1(n3085), .B0(n2828), .B1(n3087), .Y(n2877) );
  OAI22X1 U4003 ( .A0(n2832), .A1(n2839), .B0(n2836), .B1(n2831), .Y(n2881) );
  OAI22XL U4004 ( .A0(n2834), .A1(n3070), .B0(n2882), .B1(n3068), .Y(n2854) );
  OR2X1 U4005 ( .A(n2926), .B(n2925), .Y(n2902) );
  OAI22X1 U4006 ( .A0(n2929), .A1(n3177), .B0(n3179), .B1(n1045), .Y(n2909) );
  XNOR2X1 U4007 ( .A(n1038), .B(n2900), .Y(n2914) );
  OAI22XL U4008 ( .A0(n2860), .A1(n2940), .B0(n2914), .B1(n2938), .Y(n2921) );
  XNOR2X1 U4009 ( .A(n3201), .B(n3084), .Y(n2927) );
  XNOR2X1 U4010 ( .A(n1073), .B(n591), .Y(n2928) );
  NAND2X1 U4011 ( .A(n3343), .B(n3344), .Y(n2863) );
  ADDFHX1 U4012 ( .A(n2879), .B(n2878), .CI(n2877), .CO(n2876), .S(n3341) );
  XNOR2X1 U4013 ( .A(n2885), .B(n2884), .Y(n2890) );
  INVXL U4014 ( .A(n2886), .Y(n2887) );
  NAND2X1 U4015 ( .A(n2888), .B(n2887), .Y(n2889) );
  XNOR2X1 U4016 ( .A(n2897), .B(n2896), .Y(n2898) );
  BUFX2 U4017 ( .A(n2898), .Y(n3258) );
  INVXL U4018 ( .A(n2936), .Y(n2899) );
  OAI2BB1X2 U4019 ( .A0N(n3261), .A1N(n3259), .B0(n2899), .Y(n2932) );
  XNOR2X1 U4020 ( .A(n3054), .B(n2979), .Y(n2915) );
  INVXL U4021 ( .A(n3347), .Y(n2906) );
  OAI22X1 U4022 ( .A0(n3089), .A1(n3182), .B0(n3184), .B1(n2913), .Y(n3145) );
  XNOR2X1 U4023 ( .A(n3251), .B(n2900), .Y(n2941) );
  ADDFHX1 U4024 ( .A(n2924), .B(n2923), .CI(n2922), .CO(n2874), .S(n3360) );
  XNOR2X1 U4025 ( .A(n2926), .B(n2925), .Y(n3148) );
  OAI22X1 U4026 ( .A0(n2927), .A1(n3087), .B0(n3088), .B1(n3085), .Y(n3147) );
  XNOR2X1 U4027 ( .A(n2976), .B(n3173), .Y(n3066) );
  OAI22X1 U4028 ( .A0(n3066), .A1(n3177), .B0(n2929), .B1(n3179), .Y(n3133) );
  OAI22X1 U4029 ( .A0(n3071), .A1(n3068), .B0(n2931), .B1(n3070), .Y(n3131) );
  ADDFHX1 U4030 ( .A(n2933), .B(n2932), .CI(n2935), .CO(n2916), .S(n3124) );
  OAI22X1 U4031 ( .A0(n3052), .A1(n3259), .B0(n3261), .B1(n2936), .Y(n3072) );
  NOR2BX2 U4032 ( .AN(n3270), .B(n2940), .Y(n3032) );
  XNOR2X1 U4033 ( .A(n3270), .B(n2900), .Y(n2939) );
  OAI22X1 U4034 ( .A0(n2941), .A1(n2940), .B0(n2939), .B1(n2938), .Y(n3078) );
  ADDFHX4 U4035 ( .A(n2946), .B(n2947), .CI(n2945), .CO(n2949), .S(n3374) );
  ADDFHX4 U4036 ( .A(n2961), .B(n2960), .CI(n2959), .CO(n3417), .S(n3415) );
  ADDFHX4 U4037 ( .A(n2964), .B(n2963), .CI(n2962), .CO(n3421), .S(n3419) );
  OAI22X1 U4038 ( .A0(n2967), .A1(n3106), .B0(n2983), .B1(n3109), .Y(n3022) );
  XNOR2X1 U4039 ( .A(n3164), .B(n3237), .Y(n3023) );
  XNOR2X1 U4040 ( .A(n769), .B(n3181), .Y(n2978) );
  XNOR2X1 U4041 ( .A(n580), .B(n3181), .Y(n2968) );
  OAI22XL U4042 ( .A0(n3182), .A1(n2978), .B0(n2968), .B1(n3184), .Y(n3021) );
  OAI22X1 U4043 ( .A0(n3030), .A1(n3091), .B0(n3092), .B1(n3013), .Y(n3061) );
  INVXL U4044 ( .A(n3070), .Y(n2971) );
  AND2X1 U4045 ( .A(n3270), .B(n583), .Y(n2972) );
  XNOR2X1 U4046 ( .A(n3009), .B(n2974), .Y(n2977) );
  XNOR2X1 U4047 ( .A(n949), .B(n2974), .Y(n3172) );
  OAI22XL U4048 ( .A0(n3172), .A1(n3273), .B0(n2977), .B1(n3275), .Y(n3000) );
  XNOR2X1 U4049 ( .A(n579), .B(n3173), .Y(n3017) );
  OAI22XL U4050 ( .A0(n3017), .A1(n3179), .B0(n2994), .B1(n3177), .Y(n2998) );
  OAI22X1 U4051 ( .A0(n2980), .A1(n3106), .B0(n3109), .B1(n669), .Y(n3027) );
  OAI22X1 U4052 ( .A0(n2981), .A1(n3091), .B0(n3092), .B1(n589), .Y(n3026) );
  NOR2BX1 U4053 ( .AN(n3270), .B(n3106), .Y(n2992) );
  INVXL U4054 ( .A(n3092), .Y(n2984) );
  XNOR2X1 U4055 ( .A(n3006), .B(n3028), .Y(n3012) );
  AOI2BB2X1 U4056 ( .B0(n2985), .B1(n2984), .A0N(n3012), .A1N(n3091), .Y(n2986) );
  INVX2 U4057 ( .A(n2986), .Y(n2996) );
  XNOR2X1 U4058 ( .A(n3054), .B(n594), .Y(n3165) );
  XNOR2X1 U4059 ( .A(n3250), .B(n3181), .Y(n3185) );
  OAI22XL U4060 ( .A0(n2994), .A1(n3179), .B0(n3180), .B1(n3177), .Y(n3196) );
  XNOR2X1 U4061 ( .A(n3006), .B(n2512), .Y(n3056) );
  XNOR2X1 U4062 ( .A(n3009), .B(n3258), .Y(n3053) );
  XNOR2X1 U4063 ( .A(n3010), .B(n3237), .Y(n3055) );
  OAI22X1 U4064 ( .A0(n3011), .A1(n3254), .B0(n3055), .B1(n3256), .Y(n3043) );
  XNOR2X1 U4065 ( .A(n3014), .B(n3258), .Y(n3024) );
  OAI22X1 U4066 ( .A0(n3015), .A1(n3261), .B0(n3024), .B1(n3259), .Y(n3019) );
  OAI22XL U4067 ( .A0(n3017), .A1(n3177), .B0(n3016), .B1(n3179), .Y(n3018) );
  XNOR2X1 U4068 ( .A(n580), .B(n3258), .Y(n3167) );
  ADDFHX1 U4069 ( .A(n3027), .B(n3026), .CI(n3025), .CO(n3003), .S(n3169) );
  XNOR2X1 U4070 ( .A(n3029), .B(n3028), .Y(n3093) );
  OAI22X1 U4071 ( .A0(n3030), .A1(n3092), .B0(n3093), .B1(n3091), .Y(n3104) );
  OAI2BB1X1 U4072 ( .A0N(n3275), .A1N(n3273), .B0(n3031), .Y(n3114) );
  ADDHX1 U4073 ( .A(n575), .B(n3032), .CO(n3080), .S(n3113) );
  ADDFHX4 U4074 ( .A(n3042), .B(n3041), .CI(n3040), .CO(n3076), .S(n3051) );
  ADDFHX1 U4075 ( .A(n3062), .B(n3061), .CI(n3060), .CO(n3097), .S(n3064) );
  ADDFHX1 U4076 ( .A(n3065), .B(n3064), .CI(n3063), .CO(n3094), .S(n3160) );
  ADDFHX1 U4077 ( .A(n3105), .B(n3104), .CI(n3103), .CO(n3141), .S(n3118) );
  ADDFHX1 U4078 ( .A(n3115), .B(n3114), .CI(n3113), .CO(n3149), .S(n3103) );
  ADDFHX1 U4079 ( .A(n3118), .B(n3117), .CI(n3116), .CO(n3137), .S(n3121) );
  ADDFHX1 U4080 ( .A(n3124), .B(n3123), .CI(n3122), .CO(n3364), .S(n3369) );
  ADDFHX1 U4081 ( .A(n3130), .B(n3129), .CI(n3128), .CO(n3350), .S(n3125) );
  ADDFHX1 U4082 ( .A(n3136), .B(n3135), .CI(n3134), .CO(n3348), .S(n3154) );
  ADDFHX1 U4083 ( .A(n3145), .B(n3144), .CI(n3143), .CO(n3363), .S(n3353) );
  XOR3X2 U4084 ( .A(n3383), .B(n3384), .C(n3387), .Y(n3400) );
  ADDFHX1 U4085 ( .A(n3163), .B(n3162), .CI(n3161), .CO(n3046), .S(n3192) );
  XNOR2X1 U4086 ( .A(n3164), .B(n594), .Y(n3186) );
  OAI22XL U4087 ( .A0(n3165), .A1(n3271), .B0(n3186), .B1(n3269), .Y(n3205) );
  XNOR2X1 U4088 ( .A(n725), .B(n3237), .Y(n3200) );
  XNOR2X1 U4089 ( .A(n3014), .B(n2974), .Y(n3199) );
  NAND2BXL U4090 ( .AN(n3270), .B(n3173), .Y(n3174) );
  NOR2BX1 U4091 ( .AN(n3270), .B(n3179), .Y(n3216) );
  NOR2BX1 U4092 ( .AN(n645), .B(n3184), .Y(n3215) );
  OAI22XL U4093 ( .A0(n3180), .A1(n3179), .B0(n3178), .B1(n3177), .Y(n3221) );
  OAI22XL U4094 ( .A0(n3236), .A1(n3269), .B0(n3186), .B1(n3271), .Y(n3219) );
  ADDFHX1 U4095 ( .A(n3195), .B(n3194), .CI(n3193), .CO(n3187), .S(n3212) );
  ADDFHX1 U4096 ( .A(n3198), .B(n3197), .CI(n3196), .CO(n3195), .S(n3227) );
  OAI22X1 U4097 ( .A0(n3235), .A1(n3273), .B0(n3199), .B1(n3275), .Y(n3233) );
  XNOR2X1 U4098 ( .A(n1038), .B(n3253), .Y(n3218) );
  XNOR2X1 U4099 ( .A(n3201), .B(n3258), .Y(n3217) );
  OAI22XL U4100 ( .A0(n3261), .A1(n3202), .B0(n3217), .B1(n3259), .Y(n3231) );
  NOR2X1 U4101 ( .A(n3327), .B(n3326), .Y(n3209) );
  ADDHXL U4102 ( .A(n3216), .B(n3215), .CO(n3213), .S(n3301) );
  ADDFHX1 U4103 ( .A(n3227), .B(n3226), .CI(n3225), .CO(n3211), .S(n3228) );
  OAI22XL U4104 ( .A0(n3264), .A1(n3273), .B0(n3235), .B1(n3275), .Y(n3304) );
  OAI22XL U4105 ( .A0(n3238), .A1(n3256), .B0(n3254), .B1(n590), .Y(n3247) );
  NAND2BXL U4106 ( .AN(n645), .B(n3258), .Y(n3240) );
  NOR2BX1 U4107 ( .AN(n3265), .B(n3256), .Y(n3249) );
  NOR2BX1 U4108 ( .AN(n3239), .B(n3261), .Y(n3248) );
  ADDFHX1 U4109 ( .A(n3243), .B(n3242), .CI(n3241), .CO(n3230), .S(n3313) );
  OAI22XL U4110 ( .A0(n3244), .A1(n3271), .B0(n3252), .B1(n3269), .Y(n3307) );
  ADDHXL U4111 ( .A(n3249), .B(n3248), .CO(n3245), .S(n3282) );
  OAI22XL U4112 ( .A0(n3252), .A1(n3271), .B0(n3272), .B1(n3269), .Y(n3280) );
  OAI22XL U4113 ( .A0(n3272), .A1(n3271), .B0(n3270), .B1(n3269), .Y(n3283) );
  OAI22XL U4114 ( .A0(n3276), .A1(n3275), .B0(n3273), .B1(n3239), .Y(n3277) );
  ADDFX1 U4115 ( .A(n3285), .B(n3284), .CI(n3283), .CO(n3287), .S(n3278) );
  INVXL U4116 ( .A(n3286), .Y(n3290) );
  NAND2XL U4117 ( .A(n3292), .B(n3291), .Y(n3293) );
  OAI21X1 U4118 ( .A0(n3295), .A1(n3294), .B0(n3293), .Y(n3312) );
  ADDFX1 U4119 ( .A(n3304), .B(n3303), .CI(n3302), .CO(n3314), .S(n3316) );
  ADDFX1 U4120 ( .A(n3307), .B(n3306), .CI(n3305), .CO(n3308), .S(n3292) );
  NAND2XL U4121 ( .A(n3319), .B(n3320), .Y(n3906) );
  NAND2X1 U4122 ( .A(n3321), .B(n3322), .Y(n4291) );
  XNOR3X2 U4123 ( .A(n3347), .B(n3345), .C(n3346), .Y(n3390) );
  ADDFHX1 U4124 ( .A(n3353), .B(n3351), .CI(n3352), .CO(n3388), .S(n3384) );
  ADDFHX4 U4125 ( .A(n3363), .B(n3362), .CI(n3361), .CO(n3359), .S(n3393) );
  ADDFHX1 U4126 ( .A(n3369), .B(n3368), .CI(n3367), .CO(n3391), .S(n3402) );
  ADDFHX4 U4127 ( .A(n3376), .B(n3374), .CI(n3375), .CO(n3413), .S(n3411) );
  OAI21X1 U4128 ( .A0(n3379), .A1(n3378), .B0(n3377), .Y(n3381) );
  NAND2X1 U4129 ( .A(n3379), .B(n3378), .Y(n3380) );
  INVXL U4130 ( .A(n3383), .Y(n3382) );
  OAI2BB1X2 U4131 ( .A0N(n3387), .A1N(n3386), .B0(n3385), .Y(n3398) );
  ADDFHX4 U4132 ( .A(n3393), .B(n3392), .CI(n3391), .CO(n3406), .S(n3397) );
  OAI21X1 U4133 ( .A0(n3398), .A1(n3399), .B0(n3397), .Y(n3395) );
  NAND2X1 U4134 ( .A(n3398), .B(n3399), .Y(n3394) );
  NOR2X4 U4135 ( .A(n3396), .B(n3408), .Y(n3594) );
  XOR3X2 U4136 ( .A(n3399), .B(n3398), .C(n3397), .Y(n3404) );
  NOR2X2 U4137 ( .A(n3404), .B(n3403), .Y(n3591) );
  XOR3X2 U4138 ( .A(n3407), .B(n3406), .C(n3405), .Y(n3409) );
  NAND2X1 U4139 ( .A(n3412), .B(n3411), .Y(n4330) );
  NAND2X1 U4140 ( .A(n3424), .B(n3423), .Y(n3977) );
  NAND2XL U4141 ( .A(n3430), .B(n3429), .Y(n3468) );
  INVXL U4142 ( .A(n3468), .Y(n3431) );
  OAI21X1 U4143 ( .A0(n4462), .A1(n3433), .B0(n3432), .Y(n3434) );
  ADDFX1 U4144 ( .A(n3440), .B(n3439), .CI(n3438), .CO(n3511), .S(n3453) );
  ADDFX1 U4145 ( .A(n3444), .B(n3443), .CI(n3442), .CO(n3519), .S(n3455) );
  INVXL U4146 ( .A(n3447), .Y(n3448) );
  ADDFX1 U4147 ( .A(n3455), .B(n3454), .CI(n3453), .CO(n3509), .S(n3436) );
  NAND2X1 U4148 ( .A(n4068), .B(n4069), .Y(n3458) );
  INVX4 U4149 ( .A(n4469), .Y(n4379) );
  INVX2 U4150 ( .A(n3470), .Y(n4460) );
  NAND2X1 U4151 ( .A(n3972), .B(n4472), .Y(n3463) );
  NOR2X1 U4152 ( .A(n3463), .B(n4459), .Y(n3465) );
  INVXL U4153 ( .A(n3968), .Y(n4464) );
  INVXL U4154 ( .A(n4462), .Y(n3461) );
  AOI21XL U4155 ( .A0(n3461), .A1(n4472), .B0(n3460), .Y(n3462) );
  NAND2XL U4156 ( .A(Q[19]), .B(butt_a_real[0]), .Y(n3913) );
  OAI21XL U4157 ( .A0(n4277), .A1(n4274), .B0(n4278), .Y(n3475) );
  AOI21X1 U4158 ( .A0(n3476), .A1(n3915), .B0(n3475), .Y(n3606) );
  NAND2XL U4159 ( .A(n3608), .B(n3478), .Y(n3480) );
  OAI21XL U4160 ( .A0(n4337), .A1(n4334), .B0(n4338), .Y(n3477) );
  AOI21XL U4161 ( .A0(n3478), .A1(n3607), .B0(n3477), .Y(n3479) );
  NAND2XL U4162 ( .A(n3725), .B(n3482), .Y(n3496) );
  OAI21XL U4163 ( .A0(n3731), .A1(n3737), .B0(n3732), .Y(n3726) );
  OAI21XL U4164 ( .A0(n4388), .A1(n4384), .B0(n4389), .Y(n3481) );
  AOI21XL U4165 ( .A0(n3482), .A1(n3726), .B0(n3481), .Y(n3495) );
  OAI21XL U4166 ( .A0(n3495), .A1(n3497), .B0(n3498), .Y(n3483) );
  AOI21X1 U4167 ( .A0(n3494), .A1(n3484), .B0(n3483), .Y(n3986) );
  OAI21X1 U4168 ( .A0(n3986), .A1(n3982), .B0(n3983), .Y(n3981) );
  NAND2XL U4169 ( .A(Q[33]), .B(butt_a_real[14]), .Y(n3978) );
  NAND2XL U4170 ( .A(Q[34]), .B(butt_a_real[15]), .Y(n4447) );
  OAI21X1 U4171 ( .A0(n4450), .A1(n4446), .B0(n4447), .Y(n3493) );
  INVXL U4172 ( .A(n3490), .Y(n3486) );
  ADDFX1 U4173 ( .A(Q[36]), .B(butt_a_real[17]), .CI(n3489), .CO(n4089), .S(
        n4498) );
  INVX1 U4174 ( .A(n4527), .Y(n4091) );
  NAND2XL U4175 ( .A(n3491), .B(n3490), .Y(n3492) );
  INVX1 U4176 ( .A(n4602), .Y(n4568) );
  OAI21XL U4177 ( .A0(n3740), .A1(n3496), .B0(n3495), .Y(n3501) );
  INVXL U4178 ( .A(n3497), .Y(n3499) );
  NAND2XL U4179 ( .A(n3499), .B(n3498), .Y(n3500) );
  AOI22XL U4180 ( .A0(n4608), .A1(FFT2D_IN_I[16]), .B0(n4434), .B1(n4607), .Y(
        n3503) );
  NAND2XL U4181 ( .A(n4600), .B(FFT2D_IN_R[16]), .Y(n3502) );
  OAI211XL U4182 ( .A0(n1118), .A1(n4568), .B0(n3503), .C0(n3502), .Y(n3504)
         );
  ADDFX1 U4183 ( .A(n3511), .B(n3510), .CI(n3509), .CO(n3523), .S(n3456) );
  ADDFX1 U4184 ( .A(n3514), .B(n3513), .CI(n3512), .CO(n4075), .S(n3518) );
  OAI22X1 U4185 ( .A0(n3515), .A1(n4081), .B0(n4079), .B1(n4082), .Y(n4084) );
  ADDFX1 U4186 ( .A(n3520), .B(n3519), .CI(n3518), .CO(n4073), .S(n3510) );
  OAI211X1 U4187 ( .A0(n4503), .A1(n4234), .B0(n3525), .C0(n3524), .Y(
        D_real[16]) );
  ADDFX1 U4188 ( .A(n4652), .B(n3530), .CI(n3529), .CO(n3528), .S(n4007) );
  AOI22XL U4189 ( .A0(n4600), .A1(FFT2D_IN_I[18]), .B0(FFT2D_IN_R[18]), .B1(
        n4608), .Y(n3531) );
  OAI2BB1XL U4190 ( .A0N(n4607), .A1N(n4208), .B0(n3531), .Y(n3532) );
  AOI21XL U4191 ( .A0(n4007), .A1(n4602), .B0(n3532), .Y(n3533) );
  ADDFX1 U4192 ( .A(n3537), .B(n3536), .CI(n3535), .CO(n3550), .S(n2369) );
  ADDFX1 U4193 ( .A(n3540), .B(n3539), .CI(n3538), .CO(n3555), .S(n3544) );
  OAI22XL U4194 ( .A0(n3541), .A1(n4077), .B0(n3559), .B1(n4078), .Y(n3562) );
  ADDFX1 U4195 ( .A(n3546), .B(n3545), .CI(n3544), .CO(n3553), .S(n3536) );
  INVXL U4196 ( .A(n3582), .Y(n3552) );
  INVXL U4197 ( .A(n3584), .Y(n3551) );
  INVXL U4198 ( .A(n3559), .Y(n3560) );
  ADDFX1 U4199 ( .A(n3563), .B(n3562), .CI(n3561), .CO(n3574), .S(n3554) );
  INVXL U4200 ( .A(n3570), .Y(n3566) );
  OR2XL U4201 ( .A(n3578), .B(n3577), .Y(n3580) );
  NAND2XL U4202 ( .A(n3578), .B(n3577), .Y(n3579) );
  INVX2 U4203 ( .A(n3590), .Y(n4327) );
  INVXL U4204 ( .A(n3592), .Y(n3593) );
  AOI21X1 U4205 ( .A0(n4327), .A1(n3604), .B0(n3593), .Y(n3598) );
  XOR2X1 U4206 ( .A(n3598), .B(n3597), .Y(n4399) );
  AOI21X1 U4207 ( .A0(n4327), .A1(n3599), .B0(n4323), .Y(n3603) );
  XNOR2X1 U4208 ( .A(n4327), .B(n3605), .Y(n4308) );
  INVXL U4209 ( .A(n4596), .Y(n4541) );
  INVXL U4210 ( .A(n4335), .Y(n3609) );
  NAND2XL U4211 ( .A(n3609), .B(n4334), .Y(n3610) );
  INVXL U4212 ( .A(n3611), .Y(n3616) );
  NAND2XL U4213 ( .A(n3616), .B(n3614), .Y(n3612) );
  XNOR2XL U4214 ( .A(n3617), .B(n3612), .Y(n4312) );
  OR2XL U4215 ( .A(Q[19]), .B(butt_a_real[0]), .Y(n3613) );
  AND2XL U4216 ( .A(n3613), .B(n3913), .Y(n3918) );
  AOI22XL U4217 ( .A0(n4602), .A1(n4312), .B0(n4607), .B1(n3918), .Y(n3624) );
  INVXL U4218 ( .A(n3614), .Y(n3615) );
  AOI21XL U4219 ( .A0(n3617), .A1(n3616), .B0(n3615), .Y(n3622) );
  INVXL U4220 ( .A(n3618), .Y(n3620) );
  NAND2XL U4221 ( .A(n3620), .B(n3619), .Y(n3621) );
  NAND2XL U4222 ( .A(n4605), .B(n4393), .Y(n3623) );
  OAI211XL U4223 ( .A0(n4356), .A1(n4552), .B0(n3624), .C0(n3623), .Y(n3625)
         );
  INVXL U4224 ( .A(n4309), .Y(n3628) );
  AOI21X1 U4225 ( .A0(n614), .A1(n4310), .B0(n3628), .Y(n3632) );
  NAND2XL U4226 ( .A(n710), .B(n3630), .Y(n3631) );
  INVX2 U4227 ( .A(n3638), .Y(n4036) );
  INVXL U4228 ( .A(n3639), .Y(n3654) );
  INVXL U4229 ( .A(n3640), .Y(n3641) );
  AOI21X1 U4230 ( .A0(n4036), .A1(n3654), .B0(n3641), .Y(n3646) );
  INVXL U4231 ( .A(n3642), .Y(n3644) );
  NAND2XL U4232 ( .A(n3644), .B(n3643), .Y(n3645) );
  XOR2X1 U4233 ( .A(n3646), .B(n3645), .Y(n4615) );
  BUFX2 U4234 ( .A(n3647), .Y(n4029) );
  AOI21X1 U4235 ( .A0(n4036), .A1(n4029), .B0(n4031), .Y(n3653) );
  INVXL U4236 ( .A(n4033), .Y(n3651) );
  NAND2X1 U4237 ( .A(n3651), .B(n4032), .Y(n3652) );
  INVXL U4238 ( .A(n4052), .Y(n3659) );
  NAND2XL U4239 ( .A(n3659), .B(n4051), .Y(n3660) );
  INVXL U4240 ( .A(n3661), .Y(n3666) );
  NAND2XL U4241 ( .A(n3666), .B(n3664), .Y(n3662) );
  XNOR2XL U4242 ( .A(n3667), .B(n3662), .Y(n4542) );
  OR2XL U4243 ( .A(Q[0]), .B(butt_a_imag[0]), .Y(n3663) );
  AND2XL U4244 ( .A(n3663), .B(n3944), .Y(n3949) );
  AOI22XL U4245 ( .A0(n4602), .A1(n4542), .B0(n4607), .B1(n3949), .Y(n3674) );
  INVXL U4246 ( .A(n3664), .Y(n3665) );
  AOI21XL U4247 ( .A0(n3667), .A1(n3666), .B0(n3665), .Y(n3672) );
  INVXL U4248 ( .A(n3668), .Y(n3670) );
  NAND2XL U4249 ( .A(n3670), .B(n3669), .Y(n3671) );
  NAND2XL U4250 ( .A(n4605), .B(n4606), .Y(n3673) );
  OAI211XL U4251 ( .A0(n4569), .A1(n4552), .B0(n3674), .C0(n3673), .Y(n3675)
         );
  INVXL U4252 ( .A(n3677), .Y(n4540) );
  INVXL U4253 ( .A(n3692), .Y(n3693) );
  NAND2X1 U4254 ( .A(n3693), .B(n3687), .Y(n3694) );
  XOR2X2 U4255 ( .A(n4027), .B(n3694), .Y(n4578) );
  NAND2XL U4256 ( .A(n4600), .B(FFT2D_IN_I[8]), .Y(n3707) );
  OAI21XL U4257 ( .A0(n4045), .A1(n3700), .B0(n3701), .Y(n3699) );
  INVXL U4258 ( .A(n3695), .Y(n3697) );
  NAND2XL U4259 ( .A(n3697), .B(n3696), .Y(n3698) );
  AOI22XL U4260 ( .A0(n2071), .A1(n4604), .B0(n4603), .B1(n4605), .Y(n3706) );
  INVXL U4261 ( .A(n3700), .Y(n3702) );
  NAND2XL U4262 ( .A(n3702), .B(n3701), .Y(n3703) );
  AOI22XL U4263 ( .A0(n4602), .A1(n4580), .B0(n4607), .B1(n4542), .Y(n3705) );
  NAND2XL U4264 ( .A(n4608), .B(FFT2D_IN_R[8]), .Y(n3704) );
  NAND4XL U4265 ( .A(n3707), .B(n3706), .C(n3705), .D(n3704), .Y(n3708) );
  INVXL U4266 ( .A(n3713), .Y(n3715) );
  OAI2BB1X1 U4267 ( .A0N(n3717), .A1N(n4469), .B0(n3718), .Y(n3720) );
  INVXL U4268 ( .A(n3721), .Y(n3723) );
  XOR2X1 U4269 ( .A(n4379), .B(n3724), .Y(n4364) );
  NAND2XL U4270 ( .A(n4600), .B(FFT2D_IN_R[8]), .Y(n3744) );
  INVXL U4271 ( .A(n3725), .Y(n3728) );
  INVXL U4272 ( .A(n3729), .Y(n4386) );
  NAND2XL U4273 ( .A(n4386), .B(n4384), .Y(n3730) );
  OAI21XL U4274 ( .A0(n3740), .A1(n3736), .B0(n3737), .Y(n3735) );
  INVXL U4275 ( .A(n3731), .Y(n3733) );
  NAND2XL U4276 ( .A(n3733), .B(n3732), .Y(n3734) );
  AOI22XL U4277 ( .A0(n2071), .A1(n4479), .B0(n4451), .B1(n4605), .Y(n3743) );
  INVXL U4278 ( .A(n3736), .Y(n3738) );
  NAND2XL U4279 ( .A(n3738), .B(n3737), .Y(n3739) );
  AOI22XL U4280 ( .A0(n4602), .A1(n4366), .B0(n4607), .B1(n4312), .Y(n3742) );
  NAND2XL U4281 ( .A(n4608), .B(FFT2D_IN_I[8]), .Y(n3741) );
  NAND4XL U4282 ( .A(n3744), .B(n3743), .C(n3742), .D(n3741), .Y(n3745) );
  AOI21XL U4283 ( .A0(n4308), .A1(n4614), .B0(n3745), .Y(n3746) );
  OAI2BB1X2 U4284 ( .A0N(n4596), .A1N(n4364), .B0(n3746), .Y(n3747) );
  AOI21X1 U4285 ( .A0(n4485), .A1(n4598), .B0(n3747), .Y(n3748) );
  OAI2BB1X2 U4286 ( .A0N(n4594), .A1N(n4458), .B0(n3748), .Y(D_real[8]) );
  NAND2XL U4287 ( .A(n3762), .B(n4625), .Y(n3772) );
  NAND2XL U4288 ( .A(n3771), .B(lay_cnt[4]), .Y(n3773) );
  OAI211XL U4289 ( .A0(n3771), .A1(lay_cnt[4]), .B0(n3776), .C0(n3773), .Y(
        n3749) );
  INVXL U4290 ( .A(n3749), .Y(N1240) );
  NAND2XL U4291 ( .A(n604), .B(n605), .Y(n3751) );
  NAND3XL U4292 ( .A(sequence_cnt[1]), .B(sequence_cnt[0]), .C(sequence_cnt[2]), .Y(n3754) );
  OR2XL U4293 ( .A(n3964), .B(n3754), .Y(n3759) );
  XOR2XL U4294 ( .A(n3759), .B(sequence_cnt[3]), .Y(n3753) );
  NAND2XL U4295 ( .A(n3753), .B(n3768), .Y(n560) );
  NOR2BXL U4296 ( .AN(sequence_cnt[3]), .B(n3754), .Y(n3758) );
  NAND2XL U4297 ( .A(sequence_cnt[4]), .B(n3758), .Y(n3803) );
  NAND2XL U4298 ( .A(n3799), .B(n3803), .Y(n3770) );
  NAND2XL U4299 ( .A(n4678), .B(sequence_cnt[0]), .Y(n3756) );
  NAND2XL U4300 ( .A(n3799), .B(sequence_cnt[0]), .Y(n3765) );
  NAND2XL U4301 ( .A(n3765), .B(sequence_cnt[1]), .Y(n3755) );
  OAI211XL U4302 ( .A0(n3770), .A1(n3756), .B0(n3755), .C0(n3768), .Y(n562) );
  NAND2XL U4303 ( .A(n3964), .B(sequence_cnt[0]), .Y(n3757) );
  OAI211XL U4304 ( .A0(n3770), .A1(sequence_cnt[0]), .B0(n3757), .C0(n3768), 
        .Y(n563) );
  NAND2XL U4305 ( .A(n3759), .B(sequence_cnt[4]), .Y(n3760) );
  OAI211XL U4306 ( .A0(n3761), .A1(n3770), .B0(n3760), .C0(n3768), .Y(n559) );
  OAI21XL U4307 ( .A0(n3762), .A1(n4625), .B0(n3772), .Y(n3763) );
  AND2XL U4308 ( .A(sequence_cnt[1]), .B(sequence_cnt[0]), .Y(n3764) );
  NAND2XL U4309 ( .A(n4676), .B(n3764), .Y(n3769) );
  OR2XL U4310 ( .A(n4678), .B(n3765), .Y(n3766) );
  NAND2XL U4311 ( .A(sequence_cnt[2]), .B(n3766), .Y(n3767) );
  OAI211XL U4312 ( .A0(n3770), .A1(n3769), .B0(n3768), .C0(n3767), .Y(n561) );
  AOI211XL U4313 ( .A0(n3840), .A1(n3772), .B0(n4102), .C0(n3771), .Y(N1239)
         );
  AOI211XL U4314 ( .A0(n4640), .A1(n3773), .B0(n3810), .C0(n4102), .Y(N1241)
         );
  AND2XL U4315 ( .A(in_out_cnt[1]), .B(in_out_cnt[0]), .Y(n3775) );
  OR2XL U4316 ( .A(n4631), .B(in_out_cnt[2]), .Y(n3774) );
  NAND2XL U4317 ( .A(n3806), .B(n3812), .Y(n3781) );
  NAND2XL U4318 ( .A(n3810), .B(n4106), .Y(n3802) );
  INVXL U4319 ( .A(n3802), .Y(n3796) );
  INVXL U4320 ( .A(n3810), .Y(n3792) );
  NAND2XL U4321 ( .A(n3806), .B(n3789), .Y(n3791) );
  INVXL U4322 ( .A(n3806), .Y(n3790) );
  NAND2XL U4323 ( .A(n3799), .B(n3790), .Y(n3963) );
  OAI211XL U4324 ( .A0(n3792), .A1(n3847), .B0(n3791), .C0(n3963), .Y(n3794)
         );
  AOI21XL U4325 ( .A0(n3810), .A1(n4624), .B0(n3965), .Y(n3793) );
  INVXL U4326 ( .A(n3798), .Y(n3852) );
  AOI21XL U4327 ( .A0(n3852), .A1(n3847), .B0(n3810), .Y(n3800) );
  AOI211XL U4328 ( .A0(n3810), .A1(n618), .B0(n3800), .C0(n3799), .Y(n3801) );
  OAI31XL U4329 ( .A0(is_row), .A1(n3803), .A2(n3802), .B0(n3801), .Y(n3804)
         );
  OAI211XL U4330 ( .A0(n3808), .A1(n3812), .B0(n3852), .C0(n4624), .Y(n3809)
         );
  OAI21XL U4331 ( .A0(n3811), .A1(n3810), .B0(n3809), .Y(n3814) );
  OAI21XL U4332 ( .A0(n3821), .A1(n3840), .B0(n3828), .Y(n3820) );
  NAND2XL U4333 ( .A(n3826), .B(n4644), .Y(n3834) );
  AOI22XL U4334 ( .A0(n3820), .A1(is_row), .B0(n4621), .B1(sequence_cnt[2]), 
        .Y(n3825) );
  INVXL U4335 ( .A(n4650), .Y(n4627) );
  NAND2XL U4336 ( .A(n3826), .B(is_row), .Y(n4103) );
  NAND2XL U4337 ( .A(n3829), .B(n4623), .Y(n4641) );
  AOI21XL U4338 ( .A0(n4646), .A1(n4641), .B0(n3840), .Y(n3830) );
  INVXL U4339 ( .A(n3834), .Y(n3835) );
  INVXL U4340 ( .A(n4646), .Y(n3843) );
  AOI222XL U4341 ( .A0(n3835), .A1(n4625), .B0(lay_cnt[5]), .B1(n3843), .C0(
        sequence_cnt[0]), .C1(n4638), .Y(n3836) );
  NAND2XL U4342 ( .A(sequence_cnt[1]), .B(n4638), .Y(n3838) );
  OAI31XL U4343 ( .A0(n4624), .A1(is_row), .A2(n4147), .B0(n3838), .Y(n3842)
         );
  AOI2BB1X1 U4344 ( .A0N(n672), .A1N(n3840), .B0(n3839), .Y(n4620) );
  AOI211XL U4345 ( .A0(n3843), .A1(lay_cnt[4]), .B0(n3842), .C0(n3841), .Y(
        n3844) );
  INVXL U4346 ( .A(n3846), .Y(n3848) );
  OAI222XL U4347 ( .A0(n3852), .A1(n4640), .B0(n3848), .B1(n4677), .C0(n3847), 
        .C1(n1132), .Y(n4635) );
  AOI222XL U4348 ( .A0(n4635), .A1(is_row), .B0(n4621), .B1(sequence_cnt[3]), 
        .C0(n4625), .C1(n3853), .Y(n3850) );
  OAI22XL U4349 ( .A0(n3852), .A1(n4677), .B0(n672), .B1(n4640), .Y(n4643) );
  AOI222XL U4350 ( .A0(n4643), .A1(is_row), .B0(n4621), .B1(sequence_cnt[4]), 
        .C0(lay_cnt[0]), .C1(n3853), .Y(n3855) );
  INVXL U4351 ( .A(in_out_cnt[4]), .Y(n3854) );
  OAI22X1 U4352 ( .A0(n3897), .A1(n3861), .B0(n3866), .B1(n3860), .Y(
        FFT2D_OUT_I[8]) );
  OAI22X1 U4353 ( .A0(n3897), .A1(n3865), .B0(n3866), .B1(n3864), .Y(
        FFT2D_OUT_I[12]) );
  OAI22X1 U4354 ( .A0(n3897), .A1(n3863), .B0(n3866), .B1(n3862), .Y(
        FFT2D_OUT_I[4]) );
  OAI22X1 U4355 ( .A0(n3897), .A1(n3870), .B0(n3866), .B1(n3869), .Y(
        FFT2D_OUT_I[5]) );
  OAI22X1 U4356 ( .A0(n3897), .A1(n3872), .B0(n3866), .B1(n3871), .Y(
        FFT2D_OUT_I[6]) );
  OAI22X1 U4357 ( .A0(n3897), .A1(n3874), .B0(n3866), .B1(n3873), .Y(
        FFT2D_OUT_I[7]) );
  OAI22X1 U4358 ( .A0(n3897), .A1(n3878), .B0(n3866), .B1(n3877), .Y(
        FFT2D_OUT_I[9]) );
  OAI22X1 U4359 ( .A0(n3897), .A1(n3880), .B0(n3866), .B1(n3879), .Y(
        FFT2D_OUT_I[13]) );
  OAI22X1 U4360 ( .A0(n3897), .A1(n3886), .B0(n3866), .B1(n3885), .Y(
        FFT2D_OUT_I[11]) );
  OAI22X1 U4361 ( .A0(n3897), .A1(n3890), .B0(n3866), .B1(n3889), .Y(
        FFT2D_OUT_I[10]) );
  OAI22X1 U4362 ( .A0(n3897), .A1(n3892), .B0(n3866), .B1(n3891), .Y(
        FFT2D_OUT_I[3]) );
  OAI22X1 U4363 ( .A0(n3897), .A1(n3894), .B0(n3866), .B1(n3893), .Y(
        FFT2D_OUT_I[1]) );
  OAI22X1 U4364 ( .A0(n3897), .A1(n3896), .B0(n3866), .B1(n3895), .Y(
        FFT2D_OUT_I[2]) );
  OAI21XL U4365 ( .A0(n4264), .A1(n3900), .B0(n3899), .Y(n3904) );
  INVXL U4366 ( .A(n4359), .Y(n3930) );
  INVXL U4367 ( .A(n3905), .Y(n3907) );
  NAND2XL U4368 ( .A(n3907), .B(n3906), .Y(n3909) );
  XOR2XL U4369 ( .A(n3909), .B(n3908), .Y(n3923) );
  AND2XL U4370 ( .A(n4608), .B(FFT2D_IN_I[0]), .Y(n3921) );
  INVXL U4371 ( .A(n3910), .Y(n3912) );
  NAND2XL U4372 ( .A(n3912), .B(n3911), .Y(n3914) );
  XOR2XL U4373 ( .A(n3914), .B(n3913), .Y(n4342) );
  INVXL U4374 ( .A(n3915), .Y(n4276) );
  INVXL U4375 ( .A(n4275), .Y(n3916) );
  NAND2XL U4376 ( .A(n3916), .B(n4274), .Y(n3917) );
  XOR2XL U4377 ( .A(n4276), .B(n3917), .Y(n4353) );
  AOI22XL U4378 ( .A0(n4602), .A1(n3918), .B0(n2071), .B1(n4353), .Y(n3919) );
  OAI2BB1XL U4379 ( .A0N(n4605), .A1N(n4342), .B0(n3919), .Y(n3920) );
  AOI211XL U4380 ( .A0(n4600), .A1(FFT2D_IN_R[0]), .B0(n3921), .C0(n3920), .Y(
        n3922) );
  XOR2X1 U4381 ( .A(n4264), .B(n3927), .Y(n4347) );
  INVX1 U4382 ( .A(n3931), .Y(n4236) );
  OAI21XL U4383 ( .A0(n4236), .A1(n3932), .B0(n713), .Y(n3935) );
  XNOR2X1 U4384 ( .A(n3935), .B(n3934), .Y(n4573) );
  INVXL U4385 ( .A(n4573), .Y(n3962) );
  INVXL U4386 ( .A(n3936), .Y(n3938) );
  NAND2XL U4387 ( .A(n3938), .B(n3937), .Y(n3940) );
  XOR2XL U4388 ( .A(n3940), .B(n3939), .Y(n3954) );
  AND2XL U4389 ( .A(n4608), .B(FFT2D_IN_R[0]), .Y(n3952) );
  INVXL U4390 ( .A(n3941), .Y(n3943) );
  NAND2XL U4391 ( .A(n3943), .B(n3942), .Y(n3945) );
  XOR2XL U4392 ( .A(n3945), .B(n3944), .Y(n4553) );
  INVXL U4393 ( .A(n4246), .Y(n3947) );
  NAND2XL U4394 ( .A(n3947), .B(n4245), .Y(n3948) );
  AOI22XL U4395 ( .A0(n4602), .A1(n3949), .B0(n2071), .B1(n4565), .Y(n3950) );
  OAI2BB1XL U4396 ( .A0N(n4605), .A1N(n4553), .B0(n3950), .Y(n3951) );
  AOI211XL U4397 ( .A0(n4600), .A1(FFT2D_IN_I[0]), .B0(n3952), .C0(n3951), .Y(
        n3953) );
  XOR2X1 U4398 ( .A(n4236), .B(n3959), .Y(n4558) );
  OAI2BB2XL U4399 ( .B0(n3965), .B1(n3964), .A0N(is_row), .A1N(n3963), .Y(n558) );
  NAND2XL U4400 ( .A(Q[4]), .B(n4145), .Y(n3966) );
  NAND2XL U4401 ( .A(n4600), .B(FFT2D_IN_R[12]), .Y(n3990) );
  NAND2XL U4402 ( .A(n3979), .B(n3978), .Y(n3980) );
  NAND2XL U4403 ( .A(n4525), .B(n2071), .Y(n3989) );
  INVXL U4404 ( .A(n3982), .Y(n3984) );
  NAND2XL U4405 ( .A(n3984), .B(n3983), .Y(n3985) );
  XOR2X1 U4406 ( .A(n3986), .B(n3985), .Y(n4452) );
  AOI22XL U4407 ( .A0(n4605), .A1(n4452), .B0(n4434), .B1(n4602), .Y(n3988) );
  AOI22XL U4408 ( .A0(n4608), .A1(FFT2D_IN_I[12]), .B0(n4607), .B1(n4366), .Y(
        n3987) );
  NAND2XL U4409 ( .A(Q[2]), .B(n4145), .Y(n3996) );
  INVXL U4410 ( .A(n4003), .Y(n4005) );
  NOR2X1 U4411 ( .A(n4220), .B(n4563), .Y(n4015) );
  INVXL U4412 ( .A(n4008), .Y(n4010) );
  NAND2XL U4413 ( .A(n4010), .B(n4009), .Y(n4011) );
  AOI22XL U4414 ( .A0(n4608), .A1(FFT2D_IN_R[17]), .B0(n4207), .B1(n4607), .Y(
        n4013) );
  OAI2BB1XL U4415 ( .A0N(FFT2D_IN_I[17]), .A1N(n4600), .B0(n4013), .Y(n4014)
         );
  AOI211X1 U4416 ( .A0(n4602), .A1(n4226), .B0(n4015), .C0(n4014), .Y(n4016)
         );
  OAI2BB1X1 U4417 ( .A0N(n4017), .A1N(n2071), .B0(n4016), .Y(n4018) );
  NAND2X1 U4418 ( .A(n4019), .B(n4596), .Y(n4020) );
  NAND2X1 U4419 ( .A(n4599), .B(n4596), .Y(n4066) );
  BUFX2 U4420 ( .A(n4025), .Y(n4026) );
  INVXL U4421 ( .A(n4029), .Y(n4030) );
  INVXL U4422 ( .A(n4031), .Y(n4034) );
  AOI22XL U4423 ( .A0(n4600), .A1(FFT2D_IN_I[11]), .B0(n4207), .B1(n2071), .Y(
        n4062) );
  OAI21XL U4424 ( .A0(n4045), .A1(n4044), .B0(n4043), .Y(n4050) );
  INVXL U4425 ( .A(n4046), .Y(n4048) );
  NAND2XL U4426 ( .A(n4048), .B(n4047), .Y(n4049) );
  AOI22XL U4427 ( .A0(n4608), .A1(FFT2D_IN_R[11]), .B0(n4221), .B1(n4605), .Y(
        n4061) );
  NAND2XL U4428 ( .A(n4601), .B(n4602), .Y(n4060) );
  INVXL U4429 ( .A(n4054), .Y(n4056) );
  NAND2XL U4430 ( .A(n4056), .B(n4055), .Y(n4057) );
  NAND2XL U4431 ( .A(n4583), .B(n4607), .Y(n4059) );
  NAND4X1 U4432 ( .A(n4067), .B(n4066), .C(n4065), .D(n4064), .Y(D_imag[11])
         );
  INVXL U4433 ( .A(n4069), .Y(n4072) );
  INVXL U4434 ( .A(n4070), .Y(n4071) );
  INVXL U4435 ( .A(n4079), .Y(n4080) );
  ADDFX1 U4436 ( .A(n4085), .B(n4084), .CI(n4083), .CO(n4515), .S(n4074) );
  INVXL U4437 ( .A(n4509), .Y(n4088) );
  NAND2X1 U4438 ( .A(n4504), .B(n4594), .Y(n4100) );
  AOI22XL U4439 ( .A0(n4608), .A1(FFT2D_IN_I[17]), .B0(n4452), .B1(n4607), .Y(
        n4092) );
  OAI2BB1XL U4440 ( .A0N(FFT2D_IN_R[17]), .A1N(n4600), .B0(n4092), .Y(n4093)
         );
  OAI21XL U4441 ( .A0(n4624), .A1(n4104), .B0(n4103), .Y(n4105) );
  NAND2XL U4442 ( .A(n4105), .B(n4625), .Y(n4108) );
  AOI22XL U4443 ( .A0(n4106), .A1(n4145), .B0(n4621), .B1(sequence_cnt[0]), 
        .Y(n4107) );
  OAI211XL U4444 ( .A0(n4626), .A1(n4640), .B0(n4108), .C0(n4107), .Y(n4110)
         );
  NAND2XL U4445 ( .A(Q[18]), .B(n4145), .Y(n4112) );
  NAND2XL U4446 ( .A(Q[17]), .B(n4145), .Y(n4113) );
  NAND2XL U4447 ( .A(Q[16]), .B(n4145), .Y(n4114) );
  NAND2XL U4448 ( .A(Q[15]), .B(n4145), .Y(n4115) );
  NAND2XL U4449 ( .A(Q[14]), .B(n4145), .Y(n4116) );
  NAND2XL U4450 ( .A(Q[13]), .B(n4145), .Y(n4117) );
  NAND2XL U4451 ( .A(Q[12]), .B(n4145), .Y(n4118) );
  NAND2XL U4452 ( .A(Q[11]), .B(n4145), .Y(n4119) );
  NAND2XL U4453 ( .A(Q[10]), .B(n4145), .Y(n4120) );
  OAI2BB1XL U4454 ( .A0N(butt_a_imag[10]), .A1N(n4147), .B0(n4120), .Y(n483)
         );
  NAND2XL U4455 ( .A(Q[9]), .B(n4145), .Y(n4121) );
  NAND2XL U4456 ( .A(Q[8]), .B(n4145), .Y(n4122) );
  NAND2XL U4457 ( .A(Q[7]), .B(n4145), .Y(n4123) );
  NAND2XL U4458 ( .A(Q[6]), .B(n4145), .Y(n4124) );
  OAI2BB1XL U4459 ( .A0N(butt_a_imag[6]), .A1N(n4147), .B0(n4124), .Y(n549) );
  NAND2XL U4460 ( .A(Q[5]), .B(n4145), .Y(n4125) );
  NAND2XL U4461 ( .A(Q[3]), .B(n4145), .Y(n4126) );
  NAND2XL U4462 ( .A(Q[0]), .B(n4145), .Y(n4127) );
  NAND2XL U4463 ( .A(Q[36]), .B(n4145), .Y(n4128) );
  NAND2XL U4464 ( .A(Q[35]), .B(n4145), .Y(n4129) );
  NAND2XL U4465 ( .A(Q[34]), .B(n4145), .Y(n4130) );
  NAND2XL U4466 ( .A(Q[33]), .B(n4145), .Y(n4131) );
  NAND2XL U4467 ( .A(Q[32]), .B(n4145), .Y(n4132) );
  NAND2XL U4468 ( .A(Q[31]), .B(n4145), .Y(n4133) );
  NAND2XL U4469 ( .A(Q[30]), .B(n4145), .Y(n4134) );
  NAND2XL U4470 ( .A(Q[29]), .B(n4145), .Y(n4135) );
  NAND2XL U4471 ( .A(Q[28]), .B(n4145), .Y(n4136) );
  NAND2XL U4472 ( .A(Q[27]), .B(n4145), .Y(n4137) );
  NAND2XL U4473 ( .A(Q[26]), .B(n4145), .Y(n4138) );
  NAND2XL U4474 ( .A(Q[25]), .B(n4145), .Y(n4139) );
  NAND2XL U4475 ( .A(Q[24]), .B(n4145), .Y(n4140) );
  NAND2XL U4476 ( .A(Q[23]), .B(n4145), .Y(n4141) );
  NAND2XL U4477 ( .A(Q[22]), .B(n4145), .Y(n4142) );
  NAND2XL U4478 ( .A(Q[21]), .B(n4145), .Y(n4143) );
  NAND2XL U4479 ( .A(Q[20]), .B(n4145), .Y(n4144) );
  NAND2XL U4480 ( .A(Q[19]), .B(n4145), .Y(n4146) );
  OAI2BB1XL U4481 ( .A0N(butt_a_real[0]), .A1N(n4147), .B0(n4146), .Y(n501) );
  NAND2XL U4482 ( .A(Q[37]), .B(n4184), .Y(n4148) );
  NAND2XL U4483 ( .A(Q[36]), .B(n4184), .Y(n4149) );
  NAND2XL U4484 ( .A(Q[35]), .B(n4184), .Y(n4150) );
  NAND2XL U4485 ( .A(Q[34]), .B(n4184), .Y(n4151) );
  NAND2XL U4486 ( .A(Q[33]), .B(n4184), .Y(n4152) );
  NAND2XL U4487 ( .A(Q[32]), .B(n4184), .Y(n4153) );
  NAND2XL U4488 ( .A(Q[31]), .B(n4184), .Y(n4154) );
  NAND2XL U4489 ( .A(Q[30]), .B(n4184), .Y(n4155) );
  NAND2XL U4490 ( .A(Q[29]), .B(n4184), .Y(n4156) );
  NAND2XL U4491 ( .A(Q[28]), .B(n4184), .Y(n4157) );
  NAND2XL U4492 ( .A(Q[27]), .B(n4184), .Y(n4158) );
  NAND2XL U4493 ( .A(Q[26]), .B(n4184), .Y(n4159) );
  NAND2XL U4494 ( .A(Q[25]), .B(n4184), .Y(n4160) );
  NAND2XL U4495 ( .A(Q[24]), .B(n4184), .Y(n4161) );
  NAND2XL U4496 ( .A(Q[23]), .B(n4184), .Y(n4162) );
  NAND2XL U4497 ( .A(Q[22]), .B(n4184), .Y(n4163) );
  NAND2XL U4498 ( .A(Q[21]), .B(n4184), .Y(n4164) );
  NAND2XL U4499 ( .A(Q[20]), .B(n4184), .Y(n4165) );
  NAND2XL U4500 ( .A(Q[18]), .B(n4184), .Y(n4166) );
  NAND2XL U4501 ( .A(Q[17]), .B(n4184), .Y(n4167) );
  NAND2XL U4502 ( .A(Q[16]), .B(n4184), .Y(n4168) );
  NAND2XL U4503 ( .A(Q[15]), .B(n4184), .Y(n4169) );
  NAND2XL U4504 ( .A(Q[14]), .B(n4184), .Y(n4170) );
  NAND2XL U4505 ( .A(Q[13]), .B(n4184), .Y(n4171) );
  NAND2XL U4506 ( .A(Q[12]), .B(n4184), .Y(n4172) );
  NAND2XL U4507 ( .A(Q[11]), .B(n4184), .Y(n4173) );
  NAND2XL U4508 ( .A(Q[10]), .B(n4184), .Y(n4174) );
  OAI2BB1XL U4509 ( .A0N(butt_b_imag[10]), .A1N(n4186), .B0(n4174), .Y(n484)
         );
  NAND2XL U4510 ( .A(Q[9]), .B(n4184), .Y(n4175) );
  NAND2XL U4511 ( .A(Q[8]), .B(n4184), .Y(n4176) );
  NAND2XL U4512 ( .A(Q[7]), .B(n4184), .Y(n4177) );
  NAND2XL U4513 ( .A(Q[6]), .B(n4184), .Y(n4178) );
  NAND2XL U4514 ( .A(Q[5]), .B(n4184), .Y(n4179) );
  NAND2XL U4515 ( .A(Q[4]), .B(n4184), .Y(n4180) );
  NAND2XL U4516 ( .A(Q[3]), .B(n4184), .Y(n4181) );
  NAND2XL U4517 ( .A(Q[2]), .B(n4184), .Y(n4182) );
  NAND2XL U4518 ( .A(Q[1]), .B(n4184), .Y(n4183) );
  NAND2XL U4519 ( .A(Q[0]), .B(n4184), .Y(n4185) );
  NAND2XL U4520 ( .A(n655), .B(n4598), .Y(n4196) );
  NAND2X1 U4521 ( .A(n4595), .B(n4596), .Y(n4195) );
  NAND2X1 U4522 ( .A(n4599), .B(n4594), .Y(n4194) );
  NAND2XL U4523 ( .A(n4600), .B(FFT2D_IN_I[10]), .Y(n4191) );
  NAND2XL U4524 ( .A(n4601), .B(n4605), .Y(n4190) );
  AOI22XL U4525 ( .A0(n4602), .A1(n4604), .B0(n4221), .B1(n2071), .Y(n4189) );
  AOI22XL U4526 ( .A0(n4608), .A1(FFT2D_IN_R[10]), .B0(n4607), .B1(n4187), .Y(
        n4188) );
  NAND4X1 U4527 ( .A(n4196), .B(n4195), .C(n4194), .D(n4193), .Y(D_imag[10])
         );
  NAND2XL U4528 ( .A(n4600), .B(FFT2D_IN_I[12]), .Y(n4200) );
  NAND2XL U4529 ( .A(n4208), .B(n2071), .Y(n4199) );
  AOI22XL U4530 ( .A0(n4605), .A1(n4207), .B0(n4221), .B1(n4602), .Y(n4198) );
  AOI22XL U4531 ( .A0(n4608), .A1(FFT2D_IN_R[12]), .B0(n4607), .B1(n4580), .Y(
        n4197) );
  NAND2XL U4532 ( .A(n4206), .B(n2071), .Y(n4212) );
  AOI22XL U4533 ( .A0(n4608), .A1(FFT2D_IN_R[13]), .B0(n4603), .B1(n4607), .Y(
        n4211) );
  AOI22XL U4534 ( .A0(n4600), .A1(FFT2D_IN_I[13]), .B0(n4602), .B1(n4207), .Y(
        n4210) );
  NAND2XL U4535 ( .A(n4208), .B(n4605), .Y(n4209) );
  NAND4X1 U4536 ( .A(n4217), .B(n4215), .C(n4216), .D(n4218), .Y(D_imag[13])
         );
  NAND2XL U4537 ( .A(n4219), .B(n4614), .Y(n4228) );
  AOI22XL U4538 ( .A0(n4608), .A1(FFT2D_IN_R[16]), .B0(n4221), .B1(n4607), .Y(
        n4223) );
  NAND2XL U4539 ( .A(n4600), .B(FFT2D_IN_I[16]), .Y(n4222) );
  OAI211XL U4540 ( .A0(n1124), .A1(n4568), .B0(n4223), .C0(n4222), .Y(n4224)
         );
  AOI21X1 U4541 ( .A0(n4596), .A1(n4230), .B0(n4229), .Y(n4232) );
  OAI211X1 U4542 ( .A0(n4234), .A1(n4233), .B0(n4232), .C0(n4231), .Y(
        D_imag[16]) );
  INVXL U4543 ( .A(n4237), .Y(n4239) );
  NAND2XL U4544 ( .A(n4239), .B(n4238), .Y(n4240) );
  INVXL U4545 ( .A(n4416), .Y(n4242) );
  NAND2XL U4546 ( .A(n4242), .B(n4415), .Y(n4244) );
  INVXL U4547 ( .A(n4243), .Y(n4417) );
  INVXL U4548 ( .A(n4565), .Y(n4255) );
  NAND2XL U4549 ( .A(n4608), .B(FFT2D_IN_R[1]), .Y(n4254) );
  OAI21XL U4550 ( .A0(n4247), .A1(n4246), .B0(n4245), .Y(n4252) );
  INVXL U4551 ( .A(n4248), .Y(n4250) );
  NAND2XL U4552 ( .A(n4250), .B(n4249), .Y(n4251) );
  XNOR2XL U4553 ( .A(n4252), .B(n4251), .Y(n4579) );
  AOI22XL U4554 ( .A0(n4602), .A1(n4553), .B0(n2071), .B1(n4579), .Y(n4253) );
  OAI211XL U4555 ( .A0(n4255), .A1(n4563), .B0(n4254), .C0(n4253), .Y(n4256)
         );
  AOI21XL U4556 ( .A0(n4600), .A1(FFT2D_IN_I[1]), .B0(n4256), .Y(n4257) );
  OAI21XL U4557 ( .A0(n4264), .A1(n4263), .B0(n607), .Y(n4269) );
  INVXL U4558 ( .A(n4265), .Y(n4267) );
  NAND2XL U4559 ( .A(n4267), .B(n617), .Y(n4268) );
  INVXL U4560 ( .A(n4292), .Y(n4271) );
  NAND2XL U4561 ( .A(n4271), .B(n4291), .Y(n4273) );
  INVXL U4562 ( .A(n4272), .Y(n4293) );
  INVXL U4563 ( .A(n4353), .Y(n4284) );
  NAND2XL U4564 ( .A(n4608), .B(FFT2D_IN_I[1]), .Y(n4283) );
  OAI21XL U4565 ( .A0(n4276), .A1(n4275), .B0(n4274), .Y(n4281) );
  INVXL U4566 ( .A(n4277), .Y(n4279) );
  NAND2XL U4567 ( .A(n4279), .B(n4278), .Y(n4280) );
  XNOR2XL U4568 ( .A(n4281), .B(n4280), .Y(n4365) );
  AOI22XL U4569 ( .A0(n4602), .A1(n4342), .B0(n2071), .B1(n4365), .Y(n4282) );
  OAI211XL U4570 ( .A0(n4284), .A1(n4563), .B0(n4283), .C0(n4282), .Y(n4285)
         );
  AOI21XL U4571 ( .A0(n4600), .A1(FFT2D_IN_R[1]), .B0(n4285), .Y(n4286) );
  OAI21XL U4572 ( .A0(n4293), .A1(n4292), .B0(n4291), .Y(n4298) );
  NAND2XL U4573 ( .A(n4296), .B(n4295), .Y(n4297) );
  INVXL U4574 ( .A(n4365), .Y(n4301) );
  NAND2XL U4575 ( .A(n4608), .B(FFT2D_IN_I[2]), .Y(n4300) );
  AOI22XL U4576 ( .A0(n4602), .A1(n4353), .B0(n2071), .B1(n4312), .Y(n4299) );
  OAI211XL U4577 ( .A0(n4301), .A1(n4563), .B0(n4300), .C0(n4299), .Y(n4302)
         );
  AOI21XL U4578 ( .A0(n4600), .A1(FFT2D_IN_R[2]), .B0(n4302), .Y(n4303) );
  AOI22XL U4579 ( .A0(n4605), .A1(n4312), .B0(n4602), .B1(n4365), .Y(n4313) );
  OAI2BB1XL U4580 ( .A0N(n2071), .A1N(n4393), .B0(n4313), .Y(n4314) );
  OAI211XL U4581 ( .A0(n4321), .A1(n4592), .B0(n4320), .C0(n4319), .Y(
        D_real[3]) );
  INVXL U4582 ( .A(n3599), .Y(n4322) );
  INVXL U4583 ( .A(n4323), .Y(n4325) );
  AOI21X1 U4584 ( .A0(n4328), .A1(n4327), .B0(n4326), .Y(n4333) );
  INVXL U4585 ( .A(n4337), .Y(n4339) );
  NAND2XL U4586 ( .A(n4339), .B(n4338), .Y(n4340) );
  NAND2XL U4587 ( .A(n4608), .B(FFT2D_IN_I[5]), .Y(n4344) );
  AOI22XL U4588 ( .A0(n4602), .A1(n4393), .B0(n4607), .B1(n4342), .Y(n4343) );
  OAI211XL U4589 ( .A0(n4356), .A1(n4563), .B0(n4344), .C0(n4343), .Y(n4345)
         );
  NAND2XL U4590 ( .A(n4608), .B(FFT2D_IN_I[6]), .Y(n4355) );
  INVXL U4591 ( .A(n4364), .Y(n4374) );
  INVXL U4592 ( .A(n4614), .Y(n4586) );
  AOI22XL U4593 ( .A0(n4605), .A1(n4366), .B0(n4607), .B1(n4365), .Y(n4367) );
  OAI2BB1XL U4594 ( .A0N(FFT2D_IN_I[7]), .A1N(n4608), .B0(n4367), .Y(n4368) );
  AOI21XL U4595 ( .A0(n2071), .A1(n4451), .B0(n4368), .Y(n4370) );
  AOI22XL U4596 ( .A0(n4600), .A1(FFT2D_IN_R[7]), .B0(n4602), .B1(n4435), .Y(
        n4369) );
  OAI211X1 U4597 ( .A0(n1123), .A1(n4586), .B0(n4370), .C0(n4369), .Y(n4371)
         );
  INVXL U4598 ( .A(n4380), .Y(n4382) );
  NAND2XL U4599 ( .A(n4600), .B(FFT2D_IN_R[9]), .Y(n4397) );
  INVXL U4600 ( .A(n4384), .Y(n4385) );
  INVXL U4601 ( .A(n4388), .Y(n4390) );
  NAND2XL U4602 ( .A(n4390), .B(n4389), .Y(n4391) );
  NAND2XL U4603 ( .A(n4493), .B(n2071), .Y(n4396) );
  AOI22XL U4604 ( .A0(n4605), .A1(n4479), .B0(n4451), .B1(n4602), .Y(n4395) );
  AOI22XL U4605 ( .A0(n4608), .A1(FFT2D_IN_I[9]), .B0(n4607), .B1(n4393), .Y(
        n4394) );
  NAND2XL U4606 ( .A(n4600), .B(FFT2D_IN_R[10]), .Y(n4408) );
  NAND2XL U4607 ( .A(n4493), .B(n4605), .Y(n4407) );
  AOI22XL U4608 ( .A0(n4602), .A1(n4479), .B0(n4434), .B1(n2071), .Y(n4406) );
  AOI22XL U4609 ( .A0(n4608), .A1(FFT2D_IN_I[10]), .B0(n4607), .B1(n4404), .Y(
        n4405) );
  OAI21XL U4610 ( .A0(n4417), .A1(n4416), .B0(n4415), .Y(n4422) );
  INVXL U4611 ( .A(n4418), .Y(n4420) );
  NAND2XL U4612 ( .A(n4420), .B(n4419), .Y(n4421) );
  INVXL U4613 ( .A(n4579), .Y(n4425) );
  NAND2XL U4614 ( .A(n4608), .B(FFT2D_IN_R[2]), .Y(n4424) );
  AOI22XL U4615 ( .A0(n4602), .A1(n4565), .B0(n2071), .B1(n4542), .Y(n4423) );
  OAI211XL U4616 ( .A0(n4425), .A1(n4563), .B0(n4424), .C0(n4423), .Y(n4426)
         );
  AOI21XL U4617 ( .A0(n4600), .A1(FFT2D_IN_I[2]), .B0(n4426), .Y(n4427) );
  AOI22XL U4618 ( .A0(n4600), .A1(FFT2D_IN_R[11]), .B0(n4452), .B1(n2071), .Y(
        n4439) );
  AOI22XL U4619 ( .A0(n4608), .A1(FFT2D_IN_I[11]), .B0(n4434), .B1(n4605), .Y(
        n4438) );
  NAND2XL U4620 ( .A(n4493), .B(n4602), .Y(n4437) );
  NAND2XL U4621 ( .A(n4435), .B(n4607), .Y(n4436) );
  INVXL U4622 ( .A(n4446), .Y(n4448) );
  NAND2XL U4623 ( .A(n4448), .B(n4447), .Y(n4449) );
  NAND2XL U4624 ( .A(n4496), .B(n2071), .Y(n4456) );
  AOI22XL U4625 ( .A0(n4608), .A1(FFT2D_IN_I[13]), .B0(n4451), .B1(n4607), .Y(
        n4455) );
  AOI22XL U4626 ( .A0(n4600), .A1(FFT2D_IN_R[13]), .B0(n4602), .B1(n4452), .Y(
        n4454) );
  NAND2XL U4627 ( .A(n4525), .B(n4605), .Y(n4453) );
  NAND2X1 U4628 ( .A(n4472), .B(n4471), .Y(n4473) );
  AOI22XL U4629 ( .A0(n4608), .A1(FFT2D_IN_I[14]), .B0(n4479), .B1(n4607), .Y(
        n4480) );
  OAI2BB1XL U4630 ( .A0N(FFT2D_IN_R[14]), .A1N(n4600), .B0(n4480), .Y(n4481)
         );
  AOI21XL U4631 ( .A0(n4602), .A1(n4525), .B0(n4481), .Y(n4483) );
  NAND2XL U4632 ( .A(n4496), .B(n4605), .Y(n4482) );
  OAI211XL U4633 ( .A0(n1118), .A1(n4552), .B0(n4483), .C0(n4482), .Y(n4484)
         );
  AOI22XL U4634 ( .A0(n4600), .A1(FFT2D_IN_R[15]), .B0(FFT2D_IN_I[15]), .B1(
        n4608), .Y(n4492) );
  OAI2BB1XL U4635 ( .A0N(n4607), .A1N(n4493), .B0(n4492), .Y(n4494) );
  OAI211X1 U4636 ( .A0(n4503), .A1(n4502), .B0(n4501), .C0(n4500), .Y(
        D_real[15]) );
  OR2XL U4637 ( .A(n4519), .B(n4518), .Y(n4521) );
  NAND2XL U4638 ( .A(n4519), .B(n4518), .Y(n4520) );
  AOI22XL U4639 ( .A0(n4600), .A1(FFT2D_IN_R[18]), .B0(FFT2D_IN_I[18]), .B1(
        n4608), .Y(n4524) );
  OAI2BB1XL U4640 ( .A0N(n4607), .A1N(n4525), .B0(n4524), .Y(n4526) );
  AOI21XL U4641 ( .A0(n4527), .A1(n4602), .B0(n4526), .Y(n4528) );
  AOI22XL U4642 ( .A0(n4605), .A1(n4542), .B0(n4602), .B1(n4579), .Y(n4543) );
  OAI2BB1XL U4643 ( .A0N(n2071), .A1N(n4606), .B0(n4543), .Y(n4544) );
  NAND2XL U4644 ( .A(n4608), .B(FFT2D_IN_R[5]), .Y(n4555) );
  AOI22XL U4645 ( .A0(n4602), .A1(n4606), .B0(n4607), .B1(n4553), .Y(n4554) );
  NAND2XL U4646 ( .A(n4608), .B(FFT2D_IN_R[6]), .Y(n4567) );
  AOI22XL U4647 ( .A0(n4605), .A1(n4580), .B0(n4607), .B1(n4579), .Y(n4581) );
  OAI2BB1XL U4648 ( .A0N(FFT2D_IN_R[7]), .A1N(n4608), .B0(n4581), .Y(n4582) );
  AOI21XL U4649 ( .A0(n2071), .A1(n4603), .B0(n4582), .Y(n4585) );
  AOI22XL U4650 ( .A0(n4600), .A1(FFT2D_IN_I[7]), .B0(n4602), .B1(n4583), .Y(
        n4584) );
  NAND2X1 U4651 ( .A(n4595), .B(n4594), .Y(n4619) );
  NAND2XL U4652 ( .A(n4597), .B(n4596), .Y(n4618) );
  NAND2X1 U4653 ( .A(n4599), .B(n4598), .Y(n4617) );
  NAND2XL U4654 ( .A(n4600), .B(FFT2D_IN_I[9]), .Y(n4612) );
  NAND2XL U4655 ( .A(n4601), .B(n2071), .Y(n4611) );
  AOI22XL U4656 ( .A0(n4605), .A1(n4604), .B0(n4603), .B1(n4602), .Y(n4610) );
  NAND4X1 U4657 ( .A(n4619), .B(n4618), .C(n4617), .D(n4616), .Y(D_imag[9]) );
  INVXL U4658 ( .A(n4620), .Y(n4630) );
  NAND2XL U4659 ( .A(sequence_cnt[1]), .B(n4621), .Y(n4622) );
  OAI31XL U4660 ( .A0(n4624), .A1(n4623), .A2(n4677), .B0(n4622), .Y(n4629) );
  OAI22XL U4661 ( .A0(n4627), .A1(n1131), .B0(n4626), .B1(n1132), .Y(n4628) );
  OAI2BB2XL U4662 ( .B0(n4641), .B1(n1132), .A0N(sequence_cnt[3]), .A1N(n4638), 
        .Y(n4633) );
  AND2XL U4663 ( .A(n4638), .B(sequence_cnt[4]), .Y(n4639) );
  OAI2BB1XL U4664 ( .A0N(n4644), .A1N(n4643), .B0(n4642), .Y(n4645) );
  NAND2XL U4665 ( .A(n4661), .B(n4657), .Y(n4658) );
  NAND2XL U4666 ( .A(n4661), .B(n4660), .Y(n4662) );
  AOI221XL U4667 ( .A0(n4667), .A1(n4666), .B0(n4665), .B1(n4666), .C0(n4664), 
        .Y(N1166) );
endmodule

