`ifdef FUNC
`define LAT_MAX 20
`define LAT_MIN 1
`endif
`ifdef PERF
`define LAT_MAX 20
`define LAT_MIN 1
`endif

module pseudo_DRAM_data#(parameter ID_WIDTH=4, ADDR_WIDTH=32, DATA_WIDTH=16, BURST_LEN=7) (
// Glbal Signal
  	  input clk,
  	  input rst_n,
// slave interface 
      // axi write address channel 
      // src master
      input wire [ID_WIDTH-1:0]     awid_s_inf,
      input wire [ADDR_WIDTH-1:0] awaddr_s_inf,
      input wire [2:0]            awsize_s_inf,
      input wire [1:0]           awburst_s_inf,
      input wire [BURST_LEN-1:0]   awlen_s_inf,
      input wire                 awvalid_s_inf,
      // src slave
      output reg                 awready_s_inf,
      // -----------------------------
   
      // axi write data channel 
      // src master
      input wire [DATA_WIDTH-1:0]  wdata_s_inf,
      input wire                   wlast_s_inf,
      input wire                  wvalid_s_inf,
      // src slave
      output reg                  wready_s_inf,
   
      // axi write response channel 
      // src slave
      output reg  [ID_WIDTH-1:0]     bid_s_inf,
      output reg  [1:0]            bresp_s_inf,
      output reg                  bvalid_s_inf,
      // src master 
      input wire                  bready_s_inf,
      // -----------------------------
   
      // axi read address channel 
      // src master
      input wire [ID_WIDTH-1:0]     arid_s_inf,
      input wire [ADDR_WIDTH-1:0] araddr_s_inf,
      input wire [BURST_LEN-1:0]   arlen_s_inf,
      input wire [2:0]            arsize_s_inf,
      input wire [1:0]           arburst_s_inf,
      input wire                 arvalid_s_inf,
      // src slave
      output reg                 arready_s_inf,
      // -----------------------------
   
      // axi read data channel 
      // slave
      output reg [ID_WIDTH-1:0]      rid_s_inf,
      output reg [DATA_WIDTH-1:0]  rdata_s_inf,
      output reg [1:0]             rresp_s_inf,
      output reg                   rlast_s_inf,
      output reg                  rvalid_s_inf,
      // master
      input wire                  rready_s_inf
      // -----------------------------
);
// Modify your "dat" in this directory path to initialized DRAM Value

parameter DRAM_p_r = "../00_TESTBED/DRAM/DRAM_data.dat";
// Modify DRAM_R_LAT           for Initial Read Data Latency, 
//        DRAM_W_LAT           for Initial Write Data Latency
//        MAX_WAIT_READY_CYCLE for control the Upperlimit time to wait Response Ready Signal
//
//        reg [7:0] DRMA_r [0:4*64*1024-1] is the storage element in this simulation model

parameter DRAM_R_LAT = 1, DRAM_W_LAT =1, MAX_WAIT_READY_CYCLE=300;
reg	[7:0]	DRAM_r	[0:8191];   // addr from 00000000 to 0001FFF



//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
n2zmsI8cYv66xjgI32EIlELN6+7YI5WG0VDToqIiZCS7P0Neva3IUjtjU1L8MyLO
Q/R4pHhl0c7qrE1LoCtQ0AbXcUCVurMyNbZISga3ylltmvJ/Yql2ILwy1OQPA23u
UdGJ9K9vugNCc5n5KeinBPWcW98EJ4BqyUhVK/cRTMfwiB6WXFsRjs29wLtcZv3n
Qt1WG5xLsr5tpyLyP0bIQtTThg9eK8C9tuK2VLGZh/JbeShLP3RPLodCXJNliQU1
YH2mmfjO9ndL1KTv56O2z2pFCIbPeKbVnQbJGIVtHOgN3ApJN5//ahoM2bNu0NFW
Sa1MVvavvonzCDsofWaKYA==
//pragma protect end_key_block
//pragma protect digest_block
D2nlFWT4Twj9s7XJuV9E9RasT5Q=
//pragma protect end_digest_block
//pragma protect data_block
DNO8gzUIXCZc/K65iIeCKrBAUlYY4UuLnuG7yc7aUbD8aP8teFUMjlTxJq5QRPML
pEIt3hkwAMxViEb2eAcUuSt/+zpDaVDDRf+Zer0h4W1xgqTr9aIGadpIm4niz4rQ
oTNlLf4kGzPI5z4ZgsXu3Ux2LSSFXNjORy1RtcTOdhMVgedaMX/wqtQlVkFNFE7c
1qLfg2l6d/68C19EB+O3MAfyGhD0HW6EuygYwR0ED5LMnOhCa8zI7S0RFJYIAEt1
MZ46fS2V47IiGlChv3De3g8lSSxxC8ZtLPXjSEloRf4GYn+7CezfDLROFsRk/I0+
3yeqzZoLj4oamisITeH0cmoPAZBsxQkFIsdqCFx+aq3KIqeIQFsl/4N3aJBOBQEk
YUcCF9IvMEN1C2VI5LdbWtxBzPx7jGnfmZEd+m7PfSEM15aikPmDvo0fga9CV/Yp
D6G+ZfNApZXyDjUkJW4cc2A/dVbIzkaE8wJdGyXuHlBJ2W/6ZP8wmGBqyYkP4eAR
xDts0EhphnCW0vKjMWz3bYkpgJ1+8h3QcqqlFRa1J0AakAxFDwcx56V4UrUlw7iM
OO8MNiE+rQ/BW2HzbrQh8CLqbNgRX3ePABKOW7jm4JH7wVmKDrCN+5E3BGi09gop
6hzy8KR7dRmRW5K6whLwR40w3SYFts7OemN9XRjmUURc+0R1lxhcagg29OliQQrk
w/epnhuL88P3vudZpOxGHNhEf2oRC+cnw0hI7hfvAsuqFWxgSq9WZPhKVcRqtkxX
ZsLaz4daQmC+IjmP3rBL499QS6bRvUPR7M1NRJb5Yp465WjmgOm69qdB5oRCKvLB
CgZg/3nuGYuLFMln3OtMU1dqBCqMNCG0Fhd6aG2M1XNWqrmq/rWzPFjmvzFpzCec
ztxKy/xPSG33dVOmLbo5p814OZTbFP3Ps9WUDsEYo069OyDsm5lejaclSp68xgKl
4JTBm5u2H6QYr9GYB2uYeb4HtR7fOXoIq3oK8QLwPai0FjF8s98bkxMoXfkYRVr7
efVf3Cuw/UHoeepWelO/BK3LXCtIgaUVsKCn064VejdIrAqyCjGnUZmwSB3p+Qr5
KR74Xh3YzvGvcJnggCsn2o+dkP94mz+04inN6+nkqUpR8Rd/PYyNWuqdvNub39/Q
1IlLGtaxDz3qyHJtXV03zkyTVz5NSEsA1uiG1wu3TWEOr5QgERQMJxLuwn4i/ovP
Crhog3Q2eMm2ZBuwFuRSiBmwIZN0mpoIQ5XpAJ4dvefqIEnHfvrXNWhDCl19gLZL
C+/7bHtwpl71NzfEd8x+gUmm7RP0XKJphfnqTQuG+L83NPy9ImDj21pEFlX8EJru
hhZ2WXKlKsFsYD8aQujPYSIUl7ycSeCbfVGr4BW/coUaQHGpgRGpQvGmjBIB78Dz
ajUZx4ytmSfBXQfxnwKRPZGPUibwVxwUdAshauKZH7tJArPar7xM9UrZBBJycxc0
4zcNSXH3VxzbfG5C/uTtjwt6V1CCbFzVTIAJTe8Ax/YPwkBYgZn5gXcxD1p0WOe/
VY1b6fj7Oo6Q6F5mzoKRJ1NEJB5kYwDr8iSFN5Say6YK3CxGaAhLyrzOdf/zJL/T
MehHAeP+Lg3GDu8AYQiF9D7g7L7U3lXXfjj2M97OwCFgH3vGKrU1hejAON45dhoC
cW7xyDLNELBewtidMLLtaVXYNFIs5WpWbCcLNIlwn2M+3Lll71QItAuwqF7zFoGt
1dVzSJjQj3QexgFEoIXrMRgHptwUT/+JVL57eoRAtM9a1uWLU9JDTDZr3msBV0N7
TACSf3/WqgJ7Lj+FH2QEvHt+QFGysAuoRPsi+c7/ZiBbsX8Lt32AdYW6iqFQfrzI
1EcmUOeC259XNgrVy+91AkkcpIliqxrAkU9/k3tOV70jt61JDJvr7EFUudSEWNCA
PvbLRe9s18uahgpjunYEToTp4bRU1FXHWIxUbb4OMalcLlMX2jjMtUqwpZ+F9KEi
VRmtpZUD4TGSHY0+kFlUrH9lVfNRweut4pdUahf0hYg12f/GZRh/Pxw0xXr5FPGD
WtFy3YiyxRtuawNdhgb8c1nvqLupXzJJSnKmuNkfKuDMWRdQpDBeNu+QYZxrpuJx
+gwAQ907XWIi/XoVEsfh4vBYg0qpknvgsAyT2j09bxAsxz2T3NoEgbV+IFscga01
rkJIydUzB028bavkplp8GplXEoZASDspwzE3Ryr4BjnSI3NCIMZFW0PJ6LzByLbF
QUi1GMHl0wEd++wjzuiHpNLCECyc26+NAGhDIz8r2V+/ZvoBADSHXQI6ajGOC/U9
B+yQmbJvmxA489QRhQyzY6JRxDqyA0/I8uJOR6Mno04vhW3lcO54jz7HuxLamcSP
H2Vl3WWJJ/3DTUmJHc9QqC2vLAqVXb8SzzoBYztETg0isB/CVu5Dpf84E7lKKc9z
kmB7SRcYIfBCSu2uI7h+z/gZxmWe0J70D7eMWVvlo+6FxMc+OMZ81nRUCEXsVTL2
U6TPMfJexTSWm6+9HgP7m7it2gxp2xCRXlVYEKXvP05kj2oaDiMKMw2h0tNMmiGF
Ac0anlvg8zMYLC6UZ+AOoFVHmXQSmv5mhar87FoFY4QlJAa1V22RsoJgteACSzKu
Iuv2eGtR0RpdW1lEksNLYvYx+l4AD+1bJnz88aS+sHtIt9vlk/YMDVDdcEgaUOYt
8V0vO6xOjZ0SBCGbRIIiNjJK/vlercMbcal8FB6FGHlhwBQ8e/iCUW8nA/faAy/s
Kvf7LTs092fd8EWQMFSn0IGZ1qVp/m0199YqZJdqTfmEc3ssygXKVMvJiKt1VbLe
rn/LGehGKd/HDS+A4tJuFRvzbGil3Wx9uMoEq94QlrFxw1N4l6UQ1gZ/gfGQWGm5
YZunLaUJ66B9qt7i+AODG9XkigxgUbIoZ084vUZxRYyY9eFWMO6o/sbVP+P4ZO0W
OK+NvTy/86gqu9cygVd1DdJsN6KIKPdOKBFVFtLWDNEW0QprKPiHNpjgEiNunwki
catcWz1OvYQuydbHFNJSGW4BQDLdWssZxpzWmonZQbqYcbtr5WYhAqhR6hrs44Su
3ErabBuiorLZi9cmC3GQMLmvA17xUVXPae/kcw1hxZW3ADDp12VmDJJQMuenGdeD
Slyky+1azjYJt2g+uh5kq19QfBgw6XSzv8PNLqQCSFyjUdN/bCDLeCKE+z8MsCwz
Xc292zer97aN494gq+1ipiXJHThRAdoyo77dhYAFdZIsUlEBuewv7kJ897nZKZ9X
PyyaqEuPr6jzdJ1TNFTt8IfewQV6v8Uu9VtypbLOAHe3lxiVo4a/7GgMgYtabUZr
xRHYtjMyRB7FuAfs9I9uQQZlfyOx7Q5Bhov7cqoTMZMc17hqtzUm8Otbeu+h30XA
bMgbWPqob7WIuS+5E0FEpYtf96vvjomqL1WopBXPawaHMKv2wcw6FrMu3IUmytaY
4LT4uhEWPhte0uoJtOvsBGcr2LpdtHTfchb/CkuqHiLbDGbPMneNqGMK/bOiiwW0
US/Fx/Y76MvQLxjwqcvKV1MJmSmdX2VaK/zb3lUmwYcOgEoq13SQiZrkFqbPE0Td
4iOEF0OmX8qypbVqvmPneaF/EcAL3yFZNW/9+FMeF+osvF5zjwnKnV2x8I0K9cL/
y0871fvDdnp4cujHZEU+gpC02xXpiUkYe9SP7CXbtVLiU5FXxVt4d3GPd8rSBWLE
1fJIU3PpKunOa/+d/go/WwzXWlW6k5SseL9zEFW8DnXXSjumq6rTyPh9XmEUurln
gzErtbXkMWFVatxIrvKu0y7Z1vgdJfGVA8yaoGvcS/vnnqqdijaSXJPP09Vlblqp
ajxD4I8cXXlXQ+A/CoFR0XTmifkPBCZ43cd5QoOYDidgEHScZrdei+HwVh46r6L0
jSNa6yyVSSjjMckl8vNlO+h2zulzDBdpU8z/jcW7w45qZeWtUl83r8gj+Z4qXuop
FAcLq60eZNeE6OkVQpDbbgpeMJ693QW3yHhB6pPtJqygW0ridWIeePB4sK5hbdKO
pK1y9YrFqcI6M83Jxknol90swIQqSUAqB40KT4v5fSCWPxOJ8zpZ6J2Z736HJspP
73+b2X1KO+mkMsbJ3+9qBzalRCiSOfwYCGVpOYsDCi7+8mOTNMQVJhQHPgRQxqqC
EgwhTBUSi0VuY1bAx6flfCZ8bXOzUgjA9//9OkW38PbymYnCXH1VTVjIEmjz5uv3
S8nhxxMFSjUNihCEs00gNAMmhxvzhrH/EWIWsuOSLaQPrdbb1jhLWw2g3QW6ScHB
tbs+gq0W1VigTZuf9vYqrEc5otdT/T62e6AjkxwYnyY6DQvy+FCIOQCsBNuyaKpd
87vLTvUf8ZnAiP42g7p7cukLUJyC7bcfZwEUX/tMNQV6qgAjQhoavOGcn38Ny5y6
ADYutROOUxhk01cdhV1fXBWR7+W+t81cirkea5dBh/oZwenC3tkAVz5MeFz7nDLE
SDCKqM8+OjKr+mIxsQgIDTp+B3NxqS42byUP/cSIdYm0g6wEtugBBD/dQL04qlDS
0b511vRo6gpFcB2bXrIbLdqFCuGv7QKn2L/c0mtNHBzMlinPJXKOxLO9cGNRvDQH
n0Ayte05aeHRB1vDcTOkeyGfdnW8cD+Ry0BJrCEloI1elgB+ypzc3QZ+gpTUxCbl
K5ypJKbJ7BVLpfQT01XlmWPrsNFJ3ztchUA9GttBIVKSF5r0ymFNdBjgwBSGUyLi
f4AC4LGVE47NIsqBIKbfl937LYn5UqPTJ7ctARoajSMaeTQP2T4pNRGOrE5+Mllx
EfgYPe4lZ1agCqHnF4EpG/ztuqxFjkEnPu8J//sKOOXhllMMiqupndQzxcLdIUrC
O/oX0nTZxcrS6o6466yt5iQoJcT2hLFcEiW30JhcG79kl6NGPRvUgCFEVa6vUxat
Ralmk0Rog53mXPcaZXU+e6FXXNnNa0Dh2suDT1Az/MnorHElJGeMzjK5Gp9an4Oy
S7prE8eisGt54VymDzm4u7xnHeN5l+BlEgNbtyN0+o3IqljDeUPZAVlaBLQQSsTR
Zbx9ieNtEYnhWkODE7TDM/XsrfDE6fKJx4fr1oX7Mzo1QIZJV76PPtu3mZnCqdrQ
QZckv87yttTmpCYhTq7CQMgZXk77mU5F3iX/oeqNeMRuZvlnTYSHAS6kdb2k7N11
kMQWYhZG8G0qX/oKqAZuWs4tCkFn78TYYPNP8e4UjGbcSebf7V9791K4gb9e9Yvp
Vi6lXyhmac5UqLbBnUO4nRU5GfaQiTysyMEjZvTYWoVx2sYujKeCTjuIw7J4nNwi
dFfsU8jexLIzKT4jA2QieC7Z8vDCJhDlXtBDK+FwF/+l260B6xX+VGaYbpMVGBe1
xO5+jbcPeXWAdVGe5yWL3OsuybTCttDbtHyr1Y1jcUgll0jKv43Tm4K9CwApR/Qx
R1bQ9dOhOO6T/ntQk7BRxMm2w8PEI4H6wptbJkwl8bFWJzUu3x9ZqQc2U34JDrTj
xs4gc0ilJZoPHr2qc+Rlu5FdvVDVOuv7y0mxA6/pJyZSW3w3Skzc0KScPKk16nJ4
N6OxDMog+8M2S4Zq5PbcFn/AS71ZwOIVfcP6QsJZLxN+p4aNn1ItuyQU/E9RqoS9
fwA3NNTQ7RkPgTtzWLQOxCsMpmwugLQvfM2ulWAa/jHS5xcuD3WENN3XcUkgAt2S
X/yfQlPbBh1Pimu7XJOl17pbDPncGHwTb2Y1nV5MeKQgALbf5sAEcjDfhFMx1hOe
hR+pSjOACw5OgYUHHIUL+4LOqfLYUQzxx42f9VOiEefXDvpxQdzu5KYjU5GsYyXk
DGTe472nnm4fGzeGwGktnX2l+I8ASh1yJQcf692n1BJvC0Mpuwyj1zvDZM20XKPo
YzzqBXv3UaxB27Rkduvmy3BQkeLp8O0JH7m/7O8432tDt/7eABStJNslF05IWMQz
TG9OYZuodJo2cJHDbqR5Xw0Abn4hwDaC4MMengZjXugvpk/+iig2MQa/y2hmeNEx
lQCFENSy8MPgGYHYWvNSOPloBXVj8C0yZW5WyE4y0+TOAbIxXJmE1e8t6AEwlMNZ
Uiv0QANHzWVSr/W2jRu+wYwGKHrYVG33yfRACnpVCMIiS0rYoH43BICszxie47/4
XgzsKDd1cFUmrw4Dffcov7qVYQUJuSJTMX2fHRlQlqcjQnY1X1cZNR1FShHr5jZ3
OvrgYIrG8QrJVRsFfvqNInj6XreOdcHGr121iIlKb2+QYaT0VHUEpb8onEduCvXj
UthxTDx52LXH3h72IpHibhNVE+NoWDhEcGdxywHg7EKum/Q9sAdoML6MA9Ozthyg
VrrRp0oRCyEMAvjZCBcYL4PyRjqx7MQQwUl9P1Ovu74YTGJeC0f3sOrwUksuQYsQ
wC2s39WnCoYpxnwxxcNQr8Evx09FprtbEDNUbSF8OMhT0GBghDGvmedDO9be0/Cd
Yypn8JWW6XSbX3qK4C98C7NulIO4bijxure5r9TsWdrKx0zJETEygtlgL5gOfk6t
exNhj7+P/DcC2dL/xfhalo3P/jHsC4pJP8LSWH4Xb+hhGuWQL+jdzMKG8l7kvKYJ
1G+k5YqvgcNtZz4Lz706Q16jFtiKxLzUgnwLSfJtt0dbW9Ghj0WCzyQZJBEhzJxV
JdooeZQjiaDZt54gCvk76EVVvMZ/D8HBz2IzGuGLV3+TT8py0AZvq82jrvZzeM/j
hoIllDE4TF7f1SlmuJj0MWs0Hv6LP210nTz0Yx3DPLPBj2wYS4pa3oO1L7H8/vTD
4NDJtC1SCZ4ytDN+Z/hxW70f5lUACrISc4n9rI3LKuBDsDJDujDDGbMR32c3y+GG
o/AdMRXuMPPqUOWcRNJxWcnQq1I4cpM46j9rCm0Cf+D2mHTC/qSdrTRrzi75D/Y8
2cIUZ0gWMj+60BboV1bAbYPvikIEo0r4E3FETPpjRx96F+ivQ5f6lkqiRMRkoCBM
cfwr7bVsqy7OraNwoIi5kpfT7e6E0Rv1wSZHSvtYy3itdqXbsQWv26qvixkE/FYo
XNKlgYXE7e3+rK3EmXP7U4VnkJrsGG3bcDzveclq2w+WR8z12HWUNjjhnpAMUnxN
Ue0Svjjpcbp45dLCMTB3nFunCgMuOb10aRVlZYOSsqnPLaukVuEYpUY9IEw8OJTo
squ6R2VjZPXd+KsSLA/Nm5UywjciByA+qtw9ma1bYZtBVnBfEAJOF1jYF2MARZ9o
/0IXJKGSwIREj6G/LjrPkUX6I+WUEKSrlOSu+PpirV87k5pj0TYi7TiehOVks3ia
Np4kJFQoctu5+p+qCBAbc36/fM/Cq/8LnsLlbhs4QllAN/Mx6bxflLF2u7r61C5r
/o0haqQuRlO5YsrMjmgyMbOGYylyKPU0CNx9AZpB+gCf6ekMz5bZfxVXVZQZ1Hoe
/Xk0D/hwNdLGQ+/LmEUeMWCCJU8zkAR349yo637vwXsZ6hpiEML+aajG0rEA3rgm
d2MVX4ZgUwWe1D+FdkCx8Nr/fA1eQqNlxSYKpgckMaPkgX4TjJujogX/VOU9jMN9
jKeTwldSB5qIgZCgvvs88f58wijTi3jKNxIcS/jrgfiUbLK9SX6uFcb9fFICsxNE
JN5IiSTqfEYyGNIYyealcpmARYF5nmJsL9YXmomNuNpfuTCS7ZxaQqBfrl18jawC
1Rv2boBH8tFFtgESqVxuJwImSnJ3XTvK/yD3Y/Wsnn9mcosENaGPmDf1s/KiOzOM
7Xt1FbBW9zL8AIGmk3364/DdDCx/IMKV5h4l6cnAty26UKy/zc4N8EDCmW5Bxb8c
YReDYMVB7yylSm4RbaON0l/cJNEe+Kd6dcToc2V6/l3oH1gBse5sF8isC60uw7gw
iVEey4j60JIe5r+eIEgJqt8BnnNpJHZ2v96f+jYAbO3FTruPD6baGrK+9qG0pSoF
H6E/21CX5qRY0U9HR9snz/BTP9hmVzIQyOhJ/mJD1KSX8jU+ziXDjUyxA6JLmzj/
6Jj9jI0gAbl63xFRka1c4X9e07sjGmzfqaUG1pQ0B/urJhNFLiviO6GSpucngoVO
2NEdHK0GP39eMg7xxGKpiiIOahM7ciPtqY9wVgVRS64UUY8KiB1VG0J5e3J7+jm4
t6jn4Yf7G1mbevKY4voEsDItwQiO/1PfnucCO1/F+BY7emjoXGKyav5Oizrtmtj1
BOeD3LSWWf4cy2hPTsXu5M3ruHuxcolg8rW/bhYJ5bZP9IBwOGLzyq9XyaqNZds1
8i2bXUlLC+j5xIgn2miDSk6W+BGLyb5OnW3N1BJWcGGyLuIUFVpQHDQxOxleavmm
nYMQzXvvN2/Kk8dZt3NCxpgR3CGoBOI0s2CUI5u4TgBGJCA2vfrVcbCWarhqp7yN
Ix0zu+C2fgjHr1qVkkATvQysFJ/5ZNmFRCYO1dVu+GyPS1InEthqwnRwWzK+0TO2
ucNxuzW1iRr/oWE4mp8m+1wWJZFxHonBgwjJfaS5xkQ6M2AK37rq5Uj3kOPfDlxE
5PqY+YbtGEsZAwtTqrx3GBTu5S5hv5XS6IcLGQ0sgYEaHUOI1XPGhsA5+zEqVbjA
CSzPt3Iq3HY1OgC2OcdklXOjdkevNEXW6y01LSfS5wu6q3nCBmIhCrcfXVQqWAx/
3mLtbSrg0rgZ3fzfdpaG2tgtn7m989rxiZgBYv6e5bVqoez1V5y9z5J+GoFdRfaF
DW5QZZVlvXo08iDg55CtrMmCbySzMXbiM6QmtGLRbm6SNXy/ZvwtnmF8urBDmjT0
Vua/gsqktrFP5TLQxqs15+irroPbOFHQh1LhWVcp4HOWwOj3TYa5Cm9Ho+Um4BBi
0q7knxrHecFydkmafjsb5dfmsnbFGMr7LJuJ9KlKGg9iEfvsRlogzHfARp8x7NFx
1tY5g86y5jrD1QHXLpq9XJ2kqji6QxONteEfY57vJhfm0sXvYtUpZWtBL73Z7+nr
eU5qwpK5axILOanWDsT5ssJIOQ/eYfUHQCVu504kRR+gIfCPw2BKhCzSBhuVwzIq
OFz1BZ+2zAhbWr5K3nBL7QSCkbswQilpZ+6unv9RsjyQRVJEQcPUl1RedNaHWoCK
i9UNWm3svFOhvGkv8/Cdu/lIOj7JvB5/ICPX1o7+Abbqv6e7pNOVPcyCqzjuUFEI
DVTaA1Git7PCLK8sa82R8yim0kFO7LZmqRi0hJxHr9HJJQf355OljKp4RvqNQfkK
OX/d2dgf6fXug6QFto7Z/yO20ip5m9qgFXKUA91rSIQYCzsmZkCwu7fihATUuc+D
8NiI2K8edYymp64YLderiGkRkuTnDJ+ihtIg1pattYb0OvV669bv1P3p3384hbjw
JXbNhGKzw4eteaxNsaAxy4LILHYuvm22V0FSiSzsGzFrC8myqCODpiz4cC9jjJE/
C3YQ7G0jvj902HHqjuU5/kC5Louz8iyUkLMGDIx5YI0bSpKF2UTJ1cWx66F3hkAU
//DeXE7ySY5yQN8Nxl6KWGbNZGmSv8RVPrWJE0KlSpjrhrhYvyrQpEtG6KBAu/6O
5LwDqPZDoZKDY7uFjLFMHgsFoh88b2YbHmY9KPkR7HU+1HxS89apt7NTy3+lItJy
lJqy+hDK7ZLkArK/0isG1aXDcq9landFywq+XkDLplB3sRESsZ1NXX0SDxemdjcr
ttAjcFcw0vdlDj5p7+ncL7Yr4RIFa8bxftQIM768wU+jGL8VuZsCBLX+swuO9iI8
4unER8T/35ELt8rokbCF/1qwPnO+oBkWmPi92GjQAu1AksPVBLx3OyoL8ru3AJr/
B43PjTaZfji1gSpGlT0Iw7DTzqUGdyAUXroQrpmz2HwxsPcXMo7/r+pCU/VP1xeg
Gzu6mm9SNgBVxhcQbKqSoPcWKnOO7DTQUoaf+M3YqU2FwdjRMY7HT8z1X7Q2sirW
iqvVxHI6R+S1H1LdQNg4nTtuYayJPGmNtd6HnCTvU9yQgFPfwqRPFg0VB6wt7I3c
4fPDPXhmbSEds/gA6Ri5udeW1MI/fShki0e01zYb9Gp06okqmHn7sx5B08G4hI7a
PKFd0fHZbv8qqw2iSSJb8TWlnCyNzxzWzWg1RbtFrK8MgJanyijhuGtgvRQsr/HJ
kPv5yEWQzkA3VTlDH1z9pflowYdPXExjc0bWWH7E20vEJzLwNXChvzio0q13qf94
V/Vz7jKJy2njccyqeYCzTzvoas4n/SqFpMKHNUdxpcieEvsw5sV71zKMNIk43V+1
v1cOYLO3645zBwCasjEmT0eIy+GHodckUU9lHRtMrHT8kAwHF45B9U7BDTdG8VfR
mF22Ugf5oA8uWzKqSFojC3LCsoFyt/DKEz6YKIykQVjZVLevDt8MSkhjPx/MD5GA
rfTcHt1p05XJCF5YvXJwCYwbaolkWW/4yQQ+OsE34p2xaW9zpHvj7DycQO7kSYO6
5cz31/Kbe/xC9RSn1/10fmojk3vOTLq2OaOrmzBOiELH0+SN5JvH0D5A+xO3wasC
kuktNJlXAOHHqAybI61BfEt7In1BMF1qhRVm6FGr7zR5mFfyI0IN0MwP7nLyEsyl
7YfmCgE+42Y2CUyYlURHN/9QfbDtwgg3fHmGiVSNRLuS0MhDCMuJWnjPLGlEFOTl
ea8ym2uLEm8s/yAV+DEcx4+7NiR6xrs5vtfi19iDy108qtyYMhQ2Lkrl5AWS6ztt
7otOzMDJfJ3K/Zvws4DYw5/syFKUcBKnnjzqHpJAJAEEcmb3E9zNsO69GmF/yrjQ
boBv90LPl1rP+KwdtMxmeRGNINoQFrR9OmpGGt5w3MDziymzwB0fnaD6wYP8IgeD
/YLABDCA1UVFHuWuamSHSesXHOmbFpfOwt9Qp0wWaI5xW77xuKJs34Rd9PGp92SY
y5BH8ZeLYbBjqef1YL448TkEX3smEVPflgZLHrnTZuMTnhaoGW8wd5+p43EHTUw9
yl1oLzuS7Xigj6+X4kAMRkTFhGnANmFZA5n6XbUmxGPUAxtOW8vGFHocR+RMEwwq
38mGamiMxmgsUlIfquX5P9XM4jAsOOdfZU3MMDjZCV/PuAY4Wb8668vxYqOG0UCp
ZbOsnvbaeL5q+AJfdeJQwKbtaXTGDGeptUdvDCpYTmu0vTIf/ypv8uCjjS7GJ/4T
LpMj6ZH1/JozteiItCgjZ8e62Dwypt9Mq0rI81Np3drKOoewlSC6RXaAXdKPx0MU
WG1SvFgxDAE3+uVPLv/P0K7KG2XTVTjvFJi9/+DgRCOaeO63rysimYPtohPNg9se
p8qBDSiBQDlkY6SlFg+8FL4G4GiveDGm+kk6NcF8loQu9FysytUwnO97/XU9VPm+
gYbnyQbSxKYlgB2S7G1azv2TbMnrCabApON6qbH8wNblSjrhBPfzmR0ttgyfvTkh
ymhE16lcLj6IC3T+uNOJahdCvVs9FH2/Fkzv8ihNUsSDhMMMc53upuuGJQnwbhKV
3I4aEhGknp7x4eBIFEV9mc2k0qTCRcbFdVRzQgjqLK+aeKr7TSfna3cFWbWaQIMg
GZrqcnEHNfzvHQVYQCXgjoun1LX0SEGjACkIG+Hfn4j/2fS65AP288UHOSETFbZW
0doDLyP9Z5hWjDtZuQjnzcAl6skcflCpi4gbJrW8qJseIr0OKLZLnzop13+nfp9f
5hKFHhOXHVJSMsPy5UwNMFXxJtZ0FYhtZ5rtUzXBHUdJI8raU6XDhh0q2nNGncyu
Dh0S9rzYzhkKA/npKipV0gFKVmAh24oclC7IzV7GZnCq2zaaXccWCVsEp2vt54mL
qIjRcwteXmELf8CvlIf9S+9QQqCFs5+hWsIoLnK2ejQ9KVpXO6LAiqjo1CpAGcJw
5TBAKJykwL3nOmuInBdVlXFIoDk/EYXR66KPCJE8g3kFz/Kv7HN9CYtUTybfp232
ImP6G3Pt4kSMtzlPHjI1tl2fAciebNG7+YeFGZ93ZypnGAE+JmU8bYPwoxl8sUqP
+xzNV73BuFax43dJRPPB0JRzpb0UY7cCgHh1gQZ0dVWbSr6bi68eRYf8MuSgCeTx
GIHO/9iKidAKg1YgtPVPKhEW8m5C/c4qRD+Y2zks9Uj6P14YFUYmpG2gpTFlrAo6
z2kEkTbWHhRPlB+9ysGXJ4CvYVunrbRk00Pqr7QOQcLzOaUfeRgMKy++VZVSk4bt
EEdV34KSIs3AUqWUFKjP5XqHRWipEO50ngBvfbb/XXQarwlUpVmRGCZVkHT9UP60
22HJI+BK9hre91SCtWDZYzqJ/m9OEjMYfP39IU6LvgnN5u1g/eeKcWlkhGXv56Yq
x11/bfNS90/Ny99izC1z7Ou9co9UbqBuuw/qInYWrlaGlLHGXEu7maSiS3uDBlkq
ONgKU1v56ctwEpsQC/TRvQU/vPG9zCyDdsmzUIVn6YM6TsLb3mwTjs6jEKgnDFoG
oyh8D2IcPw2pVV54/wGD8lqVSdkNEVz4DTSJoCkfDQOh0/rFMVxHtis6peME8XAZ
ixGG1zCoGC06fedUwvlKt9CIcDN/jrQGkVI17g5TBSfntDOUi2IYvl0eUsivQvik
BexFNR/pYGCFO9v0/ZweJ7VJBd5gQqvTbaheYb+zaIV9gyt8DCiqhM9W6dW932xU
ulDQmgKpDqefcGyvYMA6r0hQM4B42r0GfesuZED7cVDT4oCVaHte7nYm8ilTbQLP
egCl3BA7gDoO9ek+SvgJvmJcgfzoaCrWeGdnc05qiYPNOETbD3ogUgK/cdl0plaX
kwZ2iH7cN/KrbnZZ2k1E+iDVevXqagq5I6LKGyp0TF6jlUShYyt8z1lX22olzby3
GoiDtu0pF+YIuUnWbMJZBz9V0naj3VLK94A+Yocqoh4eAUH0OkMmRxie2Bw4QCR4
mRxxUqi1KzL3TjdPjag67Pir9h/knST/VNOk6AJVKAxkoSPUu3XGOLIkwbvj+4/x
MimsIfS8GcscwQwGY4JGTNBTR54ENKiu0sVs7LWrp+7dM0w9+rhx+9vQuwBCoeVO
7OSWIF7wB961z7CEYl4s3Ptcmp1LzqEw+ZKQOY9Gs53LzZTb9Jlhihq683SzTpiZ
f/om42DmycACnnfoxCRB+zCk46sDs7vv3J3vTpdJMfBZMr06kgh5qAZBrA+Zv3Wx
W3ZSDzzBZS3iSHGBja/szBDybB0sZd//GyI3PY7PSaJVt/Iqcc1vRYhwIz2wjfZk
/ihwZS8OAPhxzsP2xZ7Yl1vozw3dGX2vLikzFT7QW24imI1nsVGjs+3M3N50B8EV
Bi7TRAjmXpxPpj2CjmI5FBLESYO6pHtI9Ux8UpB9/3iZpjKH+6UnoSTXqEbMsczp
DYCeOH8/+oWo8rV/za4a9jqt0CwEP+qRgXWVvEXaktUUK9/kr+XmjDN9bjlDVC2a
0GROw0HDfduqJ/rNGp/pRujiKhbg5ABJZQulS2tzNQIjJ1vXSPVqTYFkadwSgJ3C
HX2suRG6bQ5GhZPV8BsZPLcyEQwwyj5CPT22HGp9TqWDOPJeHYLygZIedLS6x138
ejVKa6T7YE9/Ddd0JxamukofVsddqfGtFxuApKLVG4vG90thuVtgvatXjLzo0Kd7
UgfQ5Vx4YRZncZEeA4qaoad1AtWzqLIBSGWiLnsf7FTCfw1N+FOzGxkze3RLDGPC
JxRMgeuOQjXGfz8wzKP9Mu9B50kmqA5689oC21AVQcvmn4Ko5cGijxug2GNg1jNV
gOFtojKZ4+HrlwxtHv6L3EAlJdgKn+gTxQHKqOmITOVmaT17FSaBVGpyJjKsEjfO
1On0wWScRmzGwkwJV9SKG4kMaJWThVYVX9ySR2RTy4MXmfyMoKiLEqPlPOXQWegD
Y//ehfoZyurmAPLCRe3XJHtQnFXUzOClpuNfNrah2KCeVEnVjMOsTKxFXWlzrKtP
f9KLLmueREgxOQ3C1SJyJQGcysbqIg4AgJtF5i0jLYBZrjwBeHA8Jk3gP4TJHjg6
LEzydGAC3zJsmxsg/MCXgFvLvt6XZJM4sCfA6X/OOXVc0WQhI2HDg+g2N90CyBiY
APyhi6SJW11+UIPvUIlbQ1eGskJ+PAB6EWEmEMl4TQtXhxv0iP1Vw24lGGUo3dcb
ErcHqmkq247BxXpUgCZ9N+FIc5fr1cXCpJruWA4SsZNgSpP+XC82+ecb4Z2aj4v2
i/tF7bhb8SeqpIPX7l//0AZZZ3WyGlCzXGQ6NtTZJcE9961SLs5CmBNmkCRCYYmN
dbwEgUs0lEjIe4ViCqEadihRM3BvoHQtOi8FJBKsd/kQJZZ1zPIWs9QJ4nFdzkGW
V7UzMz9gGs3pzOWWxBvvszEZmzjN0AYRDgDhNESO4WDVNXQrCzvJTPdaRI5tblvV
iZ5hCJhhns2TSIx8lIPfKiHRxCw3NUwzCKhfUQj4C996lO3LDdGxQhaqsTSABo6u
MwVpoUahjdTOxQjkfOhUJzUn5qIPWfWLCPxBX/ogGmKQRpwc2oyaG4J0Fk+APzQq
5jOqxywegaXXvS3twnOsxpMDIWRdDMV0ySdo0rJAmUTALS+EJIMEvKcbKQ9O5lzQ
8HqmeDP3VqHxeBTigaE6Zqd/s3bpX+hnGAtEj8nwg4I2LEMs0ndWToqIGXilUcVa
xndnb7IeIoEJs3tOSGxwMA1//s8yaE/JdNnkMoeqRMCdiv/Zeq4FeOVHntzYKuAL
D0k2wdTkkv76nAZkyBizQx3bi7zIYeIVIV0+yniiYM4Uq7/C/1tpjX+93I7ds3QU
DbvtpXQry4hb2nnP7T5KYT/48to4s7/ez52tq1MLl9GjSfd8S8NngNuLU8WoNkkO
bkUX2wcoAovLriKnLic9FhidL9zbvvW2n2f+tVFoTWaPQTjQx5SyfpR3jzk2e6Qw
GLtRYWmEB79fAzDt5SU8E5eey4zPQFHx9/WqSC4rphp6F1wg7DYREB0MVkWcITTI
gD8wWE01hkFhuS9DFoSVma7EVQfEyTcRX4U/j0iBcRWTh+pSZplv2+dNeqQmqGc3
kXwUpAomIgaw2gOkB/tRFlK5TWbExJplfaKbig/MrKBEo4XRI22+e77a+BqZDsGH
bXrdNsDHriC+l35Eobaz2wXNTN1QNSYLANLMmh5BCHq3LpUBM3gR4sazi9RaEdap
NIubooSuPO3SRWpOQfkjlhmCAseIt0sFr74laIpcrMrz7bYnt6yP1ESooH+Soj8k
zFCsT5QM70FM0Z/QExtaZAP11+SCmsNvLVCQOoSQf7P8GDyuFmnnHk7AwP2TbXSS
7P+kKCq+qBQ2zPy2lJus/GiMscMqMQLYOeK8SV3QJWjOE3OEi61ctl20jSWexaKK
FiGcaTd6AOQ/8zfyGnEbYMs8jFJwXxLIE3GJX7GFhtntpKSnLTvbN1aXPAmiQRs2
RBLym7cRIkYPpTmBVVghjCrsiz8h2Nk5ah5GwRuPcbSInCz0Xqr2ApTX9dLpCeNY
HON1746FG9SkOo9lZXCpJba0g/ZcoSUlpVaZku+wTY4Pm/F73QRZy587lbKVB5oo
mZAqbYhX8ItxY0St74Yyk/iVzlqGIFbxzcT9aV/5L9qMFTQINCHKTQBGLoVIF+gd
JDCGminzv6tGfctMU1uZZFTw+41nXpM6gDmO7oRITymKZuQjxSI3xp25QABN9A48
2BIIMgLu+NNm6tCAhGUytx/fG9NKxCWwczGx6AVff4tpooKn/9r4wlAM9Pu+UdDK
sFytvHz31CRBvyVefKCvdmSy+K9HuN2nUvm5EEtiM8+7+q1Vo3p8764p5kLVFC11
ksaBsnHNBTlhJrd6WuMdSN87XKGsY5oo/Bn0PpxQolICubUMhQ0UVYddweeueXgZ
zHJwvNTGSuEkRwQyGzqroNbHMi6XYm6Bg1VMmiffA4FpVk5iKF+oNtkZFDq6C1UM
7/uY1LsI99sZmp0DAEewgTIcbYNdo8JxTMAST7caNHJ8bysZT2ckCgfaEYS3oWU8
wCrkJlhSziDnXSqSjxXnSjxZqjQei1rfTr81VpbofhHUywdFEIHI6OitRD/olLcB
Tgb/Jgb8SfsIvSMj2UVyL/FjgaVE5lIaPpDWYAfO+ZElTXQgSSHIwUyOUrPvgBT7
hWFH/h3ur+GlDFp/u4sD1NHajba8o0oyZmI49xKG19kg+AzqVPN0ZTECXhNQNn/h
OX1MXeELVlc3kedzCChdE69IrBMyKIuKe6E5SEmkQaeSrQPv0BJn8N82O8+hfU30
5phXJ9W27ZOFOEzGJdjtLNutZ6jf0nQ9nefYY8dSdDWrp78Mb33ieIfApXusaFHz
sothPj6MiufdOE4C4lbQkhhyeaCDVqTUjw/0bACOuclXAPfAomIvA9NIo7/H7L1y
37xhhQGlR9akigTf87da9jV9sDn3m6Ml0ji3JDxZbjIgu45ZrpfSC2HTcSor4X4i
7q/hjGT1RHXlhGscToSE0dV5jYeQ28WCMthGgc6oJOG+m0hW3cEIfVALMqg0k+5T
s7l+NY2IQ75eZxOMII6FhwEzZoNo0lU3MKNzSJDX6k3o4bWnv4WePGwfXBmn7WTB
LCYlkr5Velx8Pr6rxmcoaFASwIrNmpVA023UgzuPyDM024sxxr1y8fl65Y0JxCU5
MmvyyPM7cXCNW5a2YQRqm9HHCTSx8jycBBoy7bauZaTXCnBYtUe86hm0RCqqSpiH
NyB4O62n+pl5i8oD/ittrlvV3ZhOehSIBORf7kSf45UOSly1fZJqdieNX6JNCW9P
iMPJa5K6UrLw6iBvOgbQfFAmkQxUHMoQtdMbLiaJ67HsIXd7btCegnBVWkSfu/hG
jHNnIe+72/b43a9kNdQixdBdgYFe9cI2VrnmaOQbBvExddUhPg5JMClLpNoauI5X
Lws1tUVG3PNqUx8rw33vmDDDYhwo37y8dpT8YuyJAFnMYHYtlvAg67oDmp6dPVlD
QOS4vEDbGwj2PNBk3qDKTFhuWRf9F36Y+8Z61zSULZsb++VOhVEDpXDKzStwWbVV
uoy4qtdAixHDhTcX3+HqVMCLt9z6jC/uonRpvjbrWtrI2xHEN0Un3bKYzRstvwVc
LCFNP1Hp2DWNJmGjGcIGloou7cBdBirSYwi4PqohUXZLL15jydRdNVYffw2ZhM74
A3GzbHi0CNmw5py5NcBETLIAmh8rt+przoLwrQMeloqgFfVvFQO3Hq9wYlqucxUg
Z8Hw4mNUVo7Dsgz1uwWwAN5spM9Vz3NYEMVbpxCOM6prKrQzTVDOW67egiU2yTsb
MXar3j5cpuSzW7HQC2L3HSEOFRQ85h28rXJZ1B+pXAp5PJkWZrouFIh6gJ1E3Hdt
TCVCcTLfzHz2S58JmtK/PWSeFVkCeBoCKFYdf7zfbHgN/1KC4Z/74pal3yYu22le
nVQhmdSglhg4LBtNnlhSNp6JJfELfqZ4Su2yIscUoVZrhrLsHMkX68Sb0WyhaUB2
lUlw0HEQ48esohpsJz4Td67r+cS+B8JnLAegwVRb7Giv/5ahcKrTXOg3eaW24TOf
f5/9tgfoxMMqKELV2G5A+GjXHZ2s4UYAL0rkfRhp0RC8k7vjG77E/h1iPekY/jFV
g9ccesro4QbDmaVPCX2lUF+YJtKjh4XSNij38qbJux2TjdccgRnGVB16gMti50ga
GviCO3maOVz3BSIDVp067djlNgqk2KBYGgV7XIPH7PhQ6J7vuhaVjs4QITOKq/oH
YUtIBttLKSInwdSaDMxY1nLe2oy9ikWVWdMxbsNOE0WlTyYnM4W1NNhixKI1hLXg
dKbvONPhsxSINsQxGvZ57H7N3QjvQYXOg/ahhncFV0vOVqZYUGowp1RIEuSXkgkW
wKpeS2iKbVgd0UnCaf5bY9QrnNZdVx79bzH/incMMey84q6qAul0TzYyvQgV7nFT
xSihp4nwrAB065G3+3MvKPu2fCDwIZR3WIA5QPJafHbPTWwc2hWch51OH8imaSJu
U2PbA3umpE1PJllA2Xq6NIXQwbhpIPT3t1m93PvYU8ppJf8L+mgbIwaZxM35a8RJ
9ZhoYdkGEsdwzjZcLDiGFQOejFq9hQZ1+AaaDK8kkgp0X+bfDxvQMVPw9auMA3sL
+9NQMgdgUwO3PgeIeb4p2bcg3JJrE8gsWtZFeL0/cpLbwMgyhRsBHx7AL3IJGBV4
wNjesXrTkv4OQI51yVTwNmRTkC7/QesWQjkYVt5Qs0IR5lQsJxOhsc2xkZ3kdMmb
2RV1YT5iPwgctTUJtLl2kWm83lOwOhqXsUGNEQecO480Hk9D/THKkIeNcJwlRcyI
mfCo7HCeIfb/nNTi6m0+aeZVF9SRosyhM44Vzi3SS0A6BZmiw7Gtxqva+9647Kvs
eRb2S9ICiuPFk956VYZOAL6Y5uvcGCjQBwLbCh2RqHZ2aDnQ+nndwGhvHU+lQQ6H
/v8FDVtwaNZGTPEt8Eg+gfo6iXw6LDnurOXMkXxhzswlAEVNIT+ruwzx0MF9pOh5
ng+1JL4KxkiFvd5XgNHJ4c5ggn4lQRjeBUG+sDew1bos5VKppywh5JHic2CygUmZ
8xWNZ2Vi8gTUlPDCLLBTq+o12tCQzAvJPv1HOID7F+3qwgkFZNrxg7WVUvkU+wBe
VA2e00w3NPyMsL5B3PffyJvn6N2NK0gJzDAuG0Sj6pflQgFyul3VURvcxk9pM5kP
DE0lNCf63nIwxRRjQ5VBrB22co7meTqAn8hqZBdudtfrvLJ/BjpoSRIVPAkVdHQy
HqN8MnCVo8FuuyEnKY1EUqV4QDo5QqmPlJ4CfiReCQiUEbX5PoI8ZBaSccfLrpnD
TeEgfPpjESTgx1samSBOUHeTHLIE0kM002s7L66zVv9htp3Ke+s3EwBTBahj4KFE
psqvWaTBM2AP7Va9Ctj5gDYc46Ou/Bhs9I3WD3Kdn10buQi9E1N9x4YwyJ30TMQe
cQNaBrfGX1MBY0DVbVCuJeM/bYJea/pUXvOc2L85jYDIYZ60Zwh5nX+a+elF+gPs
70HXp+hOyQsKgancF2y4TPIJFyH6NSjKXcNtWztsZDa2a+J0fSvR9575fbeN1IGL
RWUVn91dKvU7aGFby6WaAEWg0700RzucnyJpG7A0t0qs/ZWP6HIOTUoqpY2W5pFW
lo8JYRAQH6LqoGOvkcj+5qwArrwonrLURj1/VavP3Q3I+FaFtppNu8X0Iw96pl59
OxR2AiVwvfgiIacH3X/cLaYz/ynzoCa5j2+c2NbK8aqUhj5wrJvyIxABMtgosona
hv45cp47k5tFvqbsLK0ULNVcdzbw9jYNPiPmIA9RHaH20F8eRUBAP3EJcmOmO9ez
9Xendxm6Z4cJl/rekL5/r4wCJhPjg9iBt3Z6GDeg1Ex0aaB21lmQtK8g9Z7Goyos
iJ13ZzSD11gUMpfBEJKjlQ3eQcA7Xy9JeY5bKh20vYAK8rk16boTMaOsZZFamoXu
YjHlNA5qrcqs37NL0JDTNv4gK3AEL0eT2JfcB74xnRKE73JDFB8tr66e/IwhpAYb
Rgk68SvBg6EyJXg+dMYgBgkCKfwwVErXjD7/4fMATOXdoIZIw3JvwjLLpCAfOWmn
BpAn1mRIwr9bVRL/JGsLlvoXWe6C2zXgallEYX/iq7Yco7JRCC5aV+cf/vhHd5qT
0Td13ik5a1q4gfz6Ff7uGuzR01DhX7VlXhPhfF6NlUQLcqQRpATTeunTGyKOr0td
yKOt6KXP5jwu3fF2wkVbzzved4pe9oG8wXrq0R2B04JdwEXDOf+9um7jJS+QL0RB
zxWlt+XQggRLXaKNWfM+PvO5je1Q5QbBsAi/FyiKV1hl26h024kcEaqHyY1hHpHN
CN0w/gTLRHnoafLfISyfJK7ECCXw6Cya0sqIWxDupZS7K8tkKwZPm63jKcE734XK
EuamOsjwcNNbCeUK6cW9C4PR19lKDG570KvH5uMnUxGuh7Ry+FSlFuy/F3zzmsln
pxxHfdevGTzFyHcM6A3c7vd9hirdSsZwTEIdzcIVZanO6Z32CSfXl+acr7dVIUF8
9Om8ryEd8aHgxGIWEoAIS+MPX7S+hmCQT0+1X8348gBfPe7nlXFN5OEl1mUnBzxW
izwg1jume5ZozqvpJQZzauql59vJLc91GBVx3Y+qzp4WVk0bOh+leatAxH5TjoDW
mjjVDOVuy4vLhKQF7xlS3TTAEQ2hxwzEuQcrptJ0qYsHg7zhFqUvElmOUL+YQ5jX
HEKydO3l7W+WcM22w9FNE+DRLuRDxYnR88jpigWIIEUS7hp3oRIrzlUCQeT2D8fv
ROMOISh/+nsRFWZGDXMKfqDHU11lRgZrDT1UWErHht6eVZNwBNDoAWVICepy1Zrz
nHgQKVVZYdh2nedgBZJmqWo9yQ2R6mNiP8evT2/rAd5jgPbEZ+UIpfHo1d5uyKlb
k75LVOdC5gNBjZzr6bCc1K/S2cFt9XQiQlrJv4Z7r9RlZ7bxCXAsSMg/1/LA4hUN
SFHvyrNgejb1XgcG7E/qOm9riM+UsIrPKapC9qbMvpTK6/WtJxlZa+sjmxw0gjQd
kodGOvgKbD+0cGku5a/pHGHeuO9lGkwAd+BnBUiZSemlQAtmdy5P2tVpsmCT7zo+
/qspMi+3MIf8EeafsxoH+S+clurVMTR2ZRgVjo9wzpGkmIVFOBzym+Tm4wO/GHn2
5rvNUZ8mGXjOprB6MMbx3yJn4HEmJXKSFMeN/YS/BgMOrynXJdsgRE8ZeYzaNW/r
QrJ56GvGRihBqxTnPTLIuhMrsyFx525d+CDxG6Uf3Sr2lhdLTeLuSpX65bb6kTb5
ItWfVSHqqvwq7/GcTQGfl1/diFrehQ0Jpdd+pqFaAt3rNK+yrGMy68eHjS5JL3yC
LeZ3+uZ2cbR8/rU+9Gh83tM5ebqz45uTKASSTD0Hby6X3K2Msltmk7e9HSztTBAq
nH2OZLAMCEue61uAr2nxE4v8XP1o1z094Bk7dvOLV/9UykcV7IE/I07phZM3xIiX
hqa4B+fjs6PhF4mp1YMQBE/UxgBkzAvyCud5O19GeZG9JW2hMMdcNUlraBmhWE1Z
G/VHb62Jdr00k5usD7XwfNG7wGWTAcIt99SFPmHRqa69AhM0DIBMMCS7CbfzQKuO
E02SBjPzGToZCeCzCEPKVgEXNokROmOl68vIdqyr+RDpAiTrUoPZVP6xSFNlVDfp
oG1sdC9ywQ6aqve8c/cT4dnQsdgWvpZPE96hfwffZlgvOZQINEEYx4Hu8DEtuO0I
gSahWzAbJAypZAEGeqMhImTwHcQ9bi0RwmcepgKAGecbTIYpET3Q3VDDwc4c4v9F
uOdvL6nd2iJO9LVGKDV0F7Fksr1jgsbACtBvy1Dd0Uxs3Rb7RMj/CzsdP2DAvGy/
9iuPQW7YucQIiiJatnKyYeGIPlpgFHG4fHdmQXbAuNVXH4i6l9RoXO2un9aIaaFu
Jpw/zL1xcvsWu29U3EmhJlTULXe3P0cjO+6aMczd7DPGsXEVpAJAyZSaOPfF7lZ+
gYJF2HE10jUAHRcOCmZ0ZTNi5VYjK7r32vsCBC4s8wiElVCl1I5a2vSk26V8WqMj
Hi4my1CD8qNMOqON0jxyy5O9KViSVUCh3dZSU4eQ2PdiwwOZ4FzTJ+fREtsWSot7
er+pk2DXYFwxAUUr9pZWPhXVWPiTNY4e8fuRTChGkbgZr+QzSQL15FTVP4TgBS91
4dpPhwHy1Wxg+tt2LOTSi5OhsSkWGCol4j8DOeyMO4zXyV743GX4sX9T2MCUiqtb
tljS+b8QepYrNEwCHiWHTw6TGYOJFxUHmwNSDvjA42ynBHnA374ILjDv/97DK8aK
SvveSac5HakfEZUglIFmKIR7Xiau4jJytCEF6/a7xNBE5xdzG5/Qwg2mCcMGg/sL
sXf7ntOuBgfcYX2mWoDXk473G41jpEw0oEljWpS+QqimgoSdkC02E4hEqlTtDFZp
G+q9LNtrKf7jPySW9X0nN2oWE0fiyB6dbM30/Amy/fCnhgZdMikVYa977xpym5Di
CCZvusSmDrohj1X6FXf8nITQnhorpp1m8clh6VXOd62Hkt0z6KkAXsH06qDFWkCW
nsnQB/ubf+ScOOB+tJCbhjIoBlSgzqR+JZ97RHay8Sa57vGdfjWRRPT40jjoATLN
aSrgc1Fx2G8Wc++ANZ8Xz5bzIbehjLUY1qB3CT7Qy6nYfCQdh7ytTe75xThdcBeZ
gA6P43E6h5Cv9WhwD0r12+KUhJMIgHpNQk+R6iQg7z23lc4mJQwMhaa8FNOasOsg
Zv84FwESl5ahTYIrPEVC3L575XDpHUls5nH7XVRwEIpjWNq4oPYzsxvlT95dZyB3
ElLbit2M2LhbkA04ypq81HcnJFIjMpMAqJxkdkDZlyRycSkkpEPSH5Qm98lznSBI
kFIc90J4r/XsiJbfmJOvMEl8IK3AtZ4IJymzG3V1Gv/d5yOT0Llh548qIH00ndy8
rmo/OahvfEdEWDSMa6/4MqcCbjluhbcq3L3GNXcKgmDP0sfqQCFEzaqJi/q5ch0e
EDjNNtOurfMp2gqHQeaQ7vn519vPaHj1SIuPSbruRFoNWVRPvbKmH3kM9QytgqFJ
V/FO2cESuqi0Pn3+ZFA0q8GBPJ7Myzg+PrIZ/sdQ8oxPeilsYf0V+7qmObKSPOnM
yhZrycNGVzT89PTgabaIiMA2usjz9zGN5ZvnxDALrQcK9guBkt9Dcdqu5F1jzEXu
FA8yPqHC6xDS5XGrsY3RIZqMC57L3RxxON9butte5iyuSKTyERaGCMd1+eoe+y24
Div975XWDPmwZwCiwr+vVkHI18Qf/FvfpogfIq8+cvRXzrDuseueN7jmlvpWXLVf
AcTEGli4OPqOGLuqThooCObh38fkqkpV+Soll6GHKzHwpjD0P2ozzRSlHIYlYmhW
bDQ+y7YRPRiRCadCTXOLtLpud1pV1cxWMWsOEiJX5Whe3WK3p7ovMACeEazKfXKx
30gjDgu5iEdVJobpJUG5NhvY+b2/B5d0yaC22VaoVR0pAZ/0DwW38zQ51XLi4nsL
wqsHGHoqdxj5Td5fU1+qw8WXWHCHofj3lWWiwOOmP3qJmNVDGr89hENm77aNvosr
JmutmSKRLmx+iDW2CUP0hAyOZd/khIENBJPzWegzehnkx7REfng43lRA4lcB7zCO
LA3wBB195X3vFKjr8Q8eBC5RlMA4yrPGD/kPdgzH5h1mKvkVKERr5eWcTKOYgRJJ
GE2dX9DHi0Sizsd0c+JKee0SodNFV+MA+V5vGqfKFrZVtWsyAuyxSxZ2kKRR6g+g
iNr3shuwkyvTkI34+C+gUt5lzRMn3KtJrfAZ9JefFFa1O5xlGMgiH46OM3TFKP3Z
Ye2XdOyxjt8FJB3pMeO+s+RnvUl1zQKwtoMIDMipvdeOyRE0pQl+kqrgUPXgxJoQ
olH4kb7/7o6HbxdXBtRqKGfDhEWM/j1Ww+b4Y2wbwBwQLUYnTr4a6AhyGGyR0yTP
FlUFMQ3OtZ2tUQv8HF0kekGL1+wIOBDDXqpyZReGW3oCB2pqwsEN7WrYkfHCPUrU
9AafacTRGrXWhg2YOO0x8Q==
//pragma protect end_data_block
//pragma protect digest_block
5PGcJTS/ghl7OMLXe2QVHrCskhM=
//pragma protect end_digest_block
//pragma protect end_protected



