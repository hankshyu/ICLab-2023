module CHIP(
  // input signals

  clk,
  rst_n,
  in_valid,
  in_valid2,
  matrix,
  matrix_size,
  i_mat_idx,
  w_mat_idx,

  // output signals

  out_valid,
  out_value 
);

input clk, rst_n;
input in_valid, in_valid2;
input matrix;
input [1:0] matrix_size;
input i_mat_idx, w_mat_idx;

output out_valid;
output out_value;

//input wires
wire C_clk, BUF_CLK;
wire C_rst_n;
wire C_in_valid, C_in_valid2;
wire C_matrix;
wire [1:0] C_matrix_size;
wire C_i_mat_idx;
wire C_w_mat_idx;
//output wires
wire C_out_valid;
wire C_out_value;


MMSA CORE(                                                                                                                                                                    
  .clk        (BUF_CLK),
  .rst_n      (C_rst_n),
  .in_valid   (C_in_valid),
  .in_valid2  (C_in_valid2),
  .matrix     (C_matrix),
  .matrix_size(C_matrix_size),
  .i_mat_idx  (C_i_mat_idx),
  .w_mat_idx  (C_w_mat_idx),

  .out_valid  (C_out_valid),
  .out_value  (C_out_value)
);

CLKBUFX20 buf0(.A(C_clk),.Y(BUF_CLK));
P8C I_CLK             ( .Y(C_clk),            .P(clk),            .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b0), .CSEN(1'b1) );
P8C I_RESET           ( .Y(C_rst_n),          .P(rst_n),          .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );

P4C I_IN_VALID        ( .Y(C_in_valid),       .P(in_valid),       .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_IN_VALID2       ( .Y(C_in_valid2),      .P(in_valid2),      .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_MATRIX          ( .Y(C_matrix),         .P(matrix),         .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_MATRIX_SIZE_0   ( .Y(C_matrix_size[0]), .P(matrix_size[0]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_MATRIX_SIZE_1   ( .Y(C_matrix_size[1]), .P(matrix_size[1]), .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_I_MAT_IDX       ( .Y(C_i_mat_idx),      .P(i_mat_idx),      .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );
P4C I_W_MAT_IDX       ( .Y(C_w_mat_idx),      .P(w_mat_idx),      .A(1'b0), .ODEN(1'b0), .OCEN(1'b0), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0) );


P8C O_OUT_VALID       ( .A(C_out_valid), 	.P(out_valid), 	 .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0));
P8C O_OUT_VALUE       ( .A(C_out_value), 	.P(out_value), 	 .ODEN(1'b1), .OCEN(1'b1), .PU(1'b1), .PD(1'b0), .CEN(1'b1), .CSEN(1'b0));

//I/O power 3.3V pads x8 (DVDD + DGND)
PVDDR VDDP0 ();
PVSSR GNDP0 ();
PVDDR VDDP1 ();
PVSSR GNDP1 ();
PVDDR VDDP2 ();
PVSSR GNDP2 ();
PVDDR VDDP3 ();
PVSSR GNDP3 ();
PVDDR VDDP4 ();
PVSSR GNDP4 ();
PVDDR VDDP5 ();
PVSSR GNDP5 ();
PVDDR VDDP6 ();
PVSSR GNDP6 ();
PVDDR VDDP7 ();
PVSSR GNDP7 ();

//Core poweri 1.8V pads x? (VDD + GND)
PVDDC VDDC0 ();
PVSSC GNDC0 ();
PVDDC VDDC1 ();
PVSSC GNDC1 ();
PVDDC VDDC2 ();
PVSSC GNDC2 ();
PVDDC VDDC3 ();
PVSSC GNDC3 ();
PVDDC VDDC4 ();
PVSSC GNDC4 ();
PVDDC VDDC5 ();
PVSSC GNDC5 ();
PVDDC VDDC6 ();
PVSSC GNDC6 ();
PVDDC VDDC7 ();
PVSSC GNDC7 ();

endmodule

/////////////////////////////////////////////////////////////
// Created by: Synopsys DC Expert(TM) in wire load mode
// Version   : T-2022.03
// Date      : Tue May  2 15:03:53 2023
/////////////////////////////////////////////////////////////


module MMSA ( clk, rst_n, in_valid, in_valid2, matrix, matrix_size, i_mat_idx, 
        w_mat_idx, out_valid, out_value );
  input [1:0] matrix_size;
  input clk, rst_n, in_valid, in_valid2, matrix, i_mat_idx, w_mat_idx;
  output out_valid, out_value;
  wire   N4522, N4523, N4524, N4525, N4526, in_slut, N4584, N4585, N4586,
         N4587, N4588, N4589, N4590, N4591, N4592, N4593, N4594, N4595, N4596,
         N4597, N4598, N4599, WEN03, WEN13, WEN23, WEN33, WEN43, WEN53, WEN63,
         WEN73, reg_invalid2_signal, N4685, N4694, N4695, N4696, N4697, N4698,
         N4699, N4700, N4701, N4702, N4778, N4779, N4780, N4781, N4782, N4783,
         N4784, N4844, N4845, N4846, N4847, N4848, N4849, N4850, N4861, N4862,
         N4863, N4864, N4865, N4866, N4867, N4878, N4879, N4880, N4881, N4882,
         N4883, N4884, N4895, N4896, N4897, N4898, N4899, N4900, N4901, N4912,
         N4913, N4914, N4915, N4916, N4917, N4918, N4929, N4930, N4931, N4932,
         N4933, N4934, N4935, N4946, N4947, N4948, N4949, N4950, N4951, N4952,
         N4963, N4964, N4965, N4966, N4967, N4968, N4969, N5006, N5008, N5010,
         N5012, N5014, N5016, N5018, N5058, N5059, N5060, N5061, N5062, N5064,
         N5067, N5068, N5069, N5070, N5071, N5072, N5075, N5076, N5077, N5078,
         N5079, N5080, N5091, N5092, N5093, N5094, N5095, N5096, N5100, N5101,
         N5102, N5103, N5104, N5107, N5108, N5109, N5110, N5111, N5112, N5118,
         N5119, N5120, N5123, N5124, N5125, N5126, N5127, N5128, N5132, N5133,
         N5134, N5135, N5136, N5139, N5140, N5141, N5142, N5143, N5144, N5145,
         N5146, N5147, N5148, N5149, N5150, N5151, N5258, N5259, N5260, N5261,
         N5262, N5263, N5264, N5265, N5266, N5267, N5268, N5269, N5270, N5271,
         N5272, N5273, N5274, N5275, N5276, N5277, N5278, N5279, N5280, N5281,
         N5282, N5283, N5284, N5285, N5286, N5287, N5288, N5289, N5290, N5291,
         N5292, N5293, N5294, N5295, N5296, N5297, N5298, N5299, N5300, N5301,
         N5302, N5303, N5304, N5305, N5306, N5307, N5308, N5309, N5310, N5311,
         N5312, N5313, N5314, N5315, N5316, N5317, N5318, N5319, N5320, N5321,
         N5322, N5323, N5324, N5325, N5326, N5327, N5328, N5329, N5330, N5331,
         N5332, N5333, N5334, N5335, N5336, N5337, N5338, N5339, N5340, N5341,
         N5342, N5343, N5344, N5345, N5346, N5347, N5348, N5349, N5350, N5351,
         N5352, N5353, N5354, N5355, N5356, N5357, N5358, N5359, N5360, N5361,
         N5362, N5363, N5364, N5365, N5366, N5367, N5368, N5369, N5370, N5371,
         N5372, N5373, N5374, N5375, N5376, N5377, N5378, N5379, N5380, N5381,
         N5382, N5383, N5384, N5385, N5387, N5388, N5389, N5390, N5391, N5392,
         N5393, N5394, N5395, N5396, N5397, N5398, N5399, N5400, N5401, N5402,
         N5420, N5421, N5422, N5423, N5424, N5425, N5426, N5427, N5428, N5429,
         N5430, N5431, N5432, N5433, N5434, N5435, N5436, N5437, N5438, N5439,
         N5440, N5441, N5442, N5443, N5444, N5445, N5446, N5447, N5448, N5449,
         N5450, N5451, N5452, N5453, N5454, N5455, N5456, N5457, N5458, N5459,
         N5461, N5462, N5463, N5464, N5465, N5466, N5467, N5468, N5469, N5470,
         N5471, N5472, N5473, N5474, N5475, N5476, N5477, N5478, N5479, N5480,
         N5481, N5482, N5483, N5484, N5485, N5486, N5487, N5488, N5489, N5490,
         N5491, N5492, N5493, N5494, N5495, N5496, N5497, N5498, N5499, N5500,
         N5502, N5503, N5504, N5505, N5506, N5507, N5508, N5509, N5510, N5511,
         N5512, N5513, N5514, N5515, N5516, N5517, N5518, N5519, N5520, N5521,
         N5522, N5523, N5524, N5525, N5526, N5527, N5528, N5529, N5530, N5531,
         N5532, N5533, N5534, N5535, N5536, N5537, N5538, N5539, N5540, N5541,
         N5683, N5684, N5685, N5686, N5687, N5688, N5689, N5690, N5691, N5692,
         N5693, N5694, N5695, N5696, N5697, N5698, N5699, N5700, N5701, N5702,
         N5703, N5704, N5705, N5706, N5707, N5708, N5709, N5710, N5711, N5712,
         N5713, N5714, N5715, N5716, N5717, N5718, N5719, N5720, N5721, N5722,
         N5724, N5725, N5726, N5727, N5728, N5729, N5730, N5731, N5732, N5733,
         N5734, N5735, N5736, N5737, N5738, N5739, N5740, N5741, N5742, N5743,
         N5744, N5745, N5746, N5747, N5748, N5749, N5750, N5751, N5752, N5753,
         N5754, N5755, N5756, N5757, N5758, N5759, N5760, N5761, N5762, N5763,
         N5765, N5766, N5767, N5768, N5769, N5770, N5771, N5772, N5773, N5774,
         N5775, N5776, N5777, N5778, N5779, N5780, N5781, N5782, N5783, N5784,
         N5785, N5786, N5787, N5788, N5789, N5790, N5791, N5792, N5793, N5794,
         N5795, N5796, N5797, N5798, N5799, N5800, N5801, N5802, N5803, N5804,
         N5806, N5807, N5808, N5809, N5810, N5811, N5812, N5813, N5814, N5815,
         N5816, N5817, N5818, N5819, N5820, N5821, N5822, N5823, N5824, N5825,
         N5826, N5827, N5828, N5829, N5830, N5831, N5832, N5833, N5834, N5835,
         N5836, N5837, N5838, N5839, N5840, N5841, N5842, N5843, N5844, N5845,
         N6171, N6172, N6173, N6174, N6175, N6176, N6177, N6178, N6179, N6180,
         N6181, N6182, N6183, N6184, N6185, N6186, N6187, N6188, N6189, N6190,
         N6191, N6192, N6193, N6194, N6195, N6196, N6197, N6198, N6199, N6200,
         N6201, N6202, N6203, N6204, N6205, N6206, N6207, N6208, N6209, N6210,
         N6212, N6213, N6214, N6215, N6216, N6217, N6218, N6219, N6220, N6221,
         N6222, N6223, N6224, N6225, N6226, N6227, N6228, N6229, N6230, N6231,
         N6232, N6233, N6234, N6235, N6236, N6237, N6238, N6239, N6240, N6241,
         N6242, N6243, N6244, N6245, N6246, N6247, N6248, N6249, N6250, N6251,
         N6253, N6254, N6255, N6256, N6257, N6258, N6259, N6260, N6261, N6262,
         N6263, N6264, N6265, N6266, N6267, N6268, N6269, N6270, N6271, N6272,
         N6273, N6274, N6275, N6276, N6277, N6278, N6279, N6280, N6281, N6282,
         N6283, N6284, N6285, N6286, N6287, N6288, N6289, N6290, N6291, N6292,
         N6294, N6295, N6296, N6297, N6298, N6299, N6300, N6301, N6302, N6303,
         N6304, N6305, N6306, N6307, N6308, N6309, N6310, N6311, N6312, N6313,
         N6314, N6315, N6316, N6317, N6318, N6319, N6320, N6321, N6322, N6323,
         N6324, N6325, N6326, N6327, N6328, N6329, N6330, N6331, N6332, N6333,
         N6335, N6336, N6337, N6338, N6339, N6340, N6341, N6342, N6343, N6344,
         N6345, N6346, N6347, N6348, N6349, N6350, N6351, N6352, N6353, N6354,
         N6355, N6356, N6357, N6358, N6359, N6360, N6361, N6362, N6363, N6364,
         N6365, N6366, N6367, N6368, N6369, N6370, N6371, N6372, N6373, N6374,
         N6376, N6377, N6378, N6379, N6380, N6381, N6382, N6383, N6384, N6385,
         N6386, N6387, N6388, N6389, N6390, N6391, N6392, N6393, N6394, N6395,
         N6396, N6397, N6398, N6399, N6400, N6401, N6402, N6403, N6404, N6405,
         N6406, N6407, N6408, N6409, N6410, N6411, N6412, N6413, N6414, N6415,
         N6417, N6418, N6419, N6420, N6421, N6422, N6423, N6424, N6425, N6426,
         N6427, N6428, N6429, N6430, N6431, N6432, N6433, N6434, N6435, N6436,
         N6437, N6438, N6439, N6440, N6441, N6442, N6443, N6444, N6445, N6446,
         N6447, N6448, N6449, N6450, N6451, N6452, N6453, N6454, N6455, N6456,
         N6458, N6459, N6460, N6461, N6462, N6463, N6464, N6465, N6466, N6467,
         N6468, N6469, N6470, N6471, N6472, N6473, N6474, N6475, N6476, N6477,
         N6478, N6479, N6480, N6481, N6482, N6483, N6484, N6485, N6486, N6487,
         N6488, N6489, N6490, N6491, N6492, N6493, N6494, N6495, N6496, N6497,
         N7419, N7429, N7430, N7431, N7432, N7433, N7434, N7475, N7476, N7477,
         N7478, N7479, N7480, N7521, N7522, N7523, N7524, N7525, N7526, N7565,
         N7566, N7567, N7568, N7569, N7570, N7606, N7607, N7608, N7609, N7610,
         N7611, N7648, N7649, N7650, N7651, N7652, N7688, N7689, N7690, N7691,
         N7692, N7693, N7727, N7728, N7729, N7730, N7731, N7764, N7765, N7766,
         N7767, N7799, N7800, N7801, N7802, N7803, N7835, N7836, N7837, N7838,
         N7839, N7840, N7871, N7872, N7873, N7874, N7875, N7907, N7908, N7909,
         N7910, N7911, N7943, N7944, N7945, N7946, N7947, N7980, N7981, N7982,
         N7983, N8480, N8517, N8518, N8519, N8520, N8521, N8522, N8523, N8524,
         N8752, N8753, N8754, N8755, N8756, N8757, N9425, N9661, N9710, N9759,
         N9808, N9857, N9906, N11045, n93, n94, n96, n98, n99, n101, n102,
         n103, n104, n107, n108, n111, n114, n115, n116, n117, n118, n119,
         n123, n132, n135, n138, n140, n141, n142, n143, n144, n164, n165,
         n166, n168, n169, n170, n171, n177, n178, n179, n180, n181, n182,
         n185, n186, n187, n188, n190, n192, n193, n194, n196, n197, n198,
         n199, n200, n202, n203, n205, n207, n210, n211, n212, n213, n214,
         n216, n219, n220, n221, n223, n224, n225, n226, n227, n229, n231,
         n239, n242, n243, n244, n245, n246, n252, n253, n260, n261, n270,
         n272, n274, n275, n276, n277, n279, n280, n282, n283, n287, n289,
         n290, n292, n293, n295, n297, n300, n301, n306, n307, n308, n309,
         n310, n313, n321, n324, n325, n326, n327, n328, n334, n335, n343,
         n344, n345, n346, n347, n349, n350, n351, n353, n354, n356, n358,
         n359, n361, n364, n365, n370, n371, n372, n373, n374, n377, n385,
         n388, n389, n390, n391, n392, n398, n399, n407, n408, n410, n411,
         n413, n415, n416, n418, n421, n422, n427, n428, n429, n430, n431,
         n434, n442, n445, n446, n447, n448, n449, n455, n456, n464, n465,
         n466, n467, n468, n470, n471, n473, n475, n476, n478, n481, n482,
         n487, n488, n489, n490, n491, n494, n502, n505, n506, n507, n508,
         n509, n515, n516, n524, n526, n527, n529, n531, n532, n534, n537,
         n538, n543, n544, n545, n546, n547, n550, n558, n561, n562, n563,
         n564, n565, n571, n572, n580, n581, n582, n583, n584, n586, n588,
         n589, n590, n591, n592, n594, n596, n597, n598, n599, n600, n601,
         n602, n604, n605, n607, n609, n610, n612, n615, n616, n621, n622,
         n623, n624, n625, n628, n636, n639, n640, n641, n642, n643, n649,
         n650, n658, n660, n661, n663, n665, n666, n668, n671, n672, n677,
         n678, n679, n680, n681, n684, n692, n695, n696, n697, n698, n699,
         n705, n706, n714, n715, n717, n718, n719, n720, n721, n722, n724,
         n725, n726, n732, n733, n734, n737, n739, n742, n743, n744, n745,
         n747, n749, n751, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n771, n772, n774,
         n775, n777, n780, n782, n784, n785, n786, n787, n788, n790, n791,
         n792, n793, n794, n797, n799, n800, n801, n802, n804, n808, n809,
         n811, n812, n814, n815, n816, n817, n818, n819, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n831, n832, n835, n836, n837,
         n838, n839, n840, n846, n849, n851, n852, n853, n854, n857, n858,
         n859, n860, n861, n862, n863, n865, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n880, n882, n883, n884,
         n888, n889, n890, n891, n895, n896, n897, n899, n900, n901, n905,
         n909, n912, n913, n917, n918, n919, n920, n921, n923, n925, n928,
         n929, n934, n1224, n1233, n1237, n1238, n1247, n1248, n1257, n1258,
         n1259, n1268, n1269, n1270, n1271, n1280, n1281, n1290, n1292, n1301,
         n1302, n1311, n1312, n1313, n1314, n1327, n1328, n1329, n1340, n1342,
         n1343, n1345, n1346, n1348, n1350, n1351, n1354, n1381, n1383, n1395,
         n1396, n1398, n1402, n1403, n1404, n1434, n1435, n1436, n1449, n1450,
         n1452, n1455, n1456, n1457, n1484, n1486, n1488, n1489, n1501, n1502,
         n1504, n1507, n1508, n1509, n1536, n1538, n1539, n1550, n1551, n1553,
         n1555, n1556, n1558, n1561, n1585, n1587, n1589, n1601, n1602, n1604,
         n1607, n1608, n1609, n1642, n1643, n1644, n1654, n1655, n1657, n1660,
         n1661, n1662, n1691, n1693, n1694, n1706, n1707, n1709, n1712, n1713,
         n1714, n1743, n1746, n1747, n1749, n1753, n1756, n1758, n1760, n1762,
         n1763, n1766, n1767, n1769, n1772, n1773, n1774, n1779, n1826, n1827,
         n1829, n1831, n1834, n1838, n1841, n1843, n1845, n1847, n1848, n1851,
         n1852, n1854, n1856, n1857, n1859, n1862, n1863, n1864, n1907, n1909,
         n1910, n1911, n1913, n1914, n1916, n1920, n1923, n1925, n1927, n1929,
         n1930, n1933, n1934, n1936, n1939, n1940, n1941, n1944, n1988, n1993,
         n1994, n1995, n1997, n2000, n2002, n2005, n2008, n2011, n2012, n2015,
         n2016, n2018, n2021, n2022, n2023, n2070, n2072, n2073, n2075, n2078,
         n2082, n2084, n2086, n2088, n2090, n2091, n2094, n2095, n2097, n2099,
         n2100, n2102, n2105, n2106, n2107, n2108, n2153, n2154, n2156, n2157,
         n2159, n2163, n2166, n2168, n2170, n2172, n2173, n2263, n2264, n2265,
         n2267, n2268, n2270, n2271, n2272, n2273, n2276, n2350, n2351, n2352,
         n2353, n2354, n2362, n2363, n2365, n2366, n2376, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2422,
         n2428, n2429, n2430, n2431, n2432, n2433, n2435, n2436, n2438, n2439,
         n2440, n2442, n2444, n2445, n2446, n2447, n2448, n2449, n2451, n2453,
         n2454, n2456, n2458, n2459, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2533, n2534, n2535, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2692, n2694, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2710, n2711, n2712, n2713, n2715, n2716, n2717, n2718, n2720, n2721,
         n2722, n2723, n2724, n2725, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2743,
         n2744, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2823, n2835, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2852,
         n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
         n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         sub_844_carry_2_, sub_844_carry_3_, sub_844_carry_4_,
         sub_844_carry_5_, sub_844_carry_6_, sub_838_carry_2_,
         sub_838_carry_3_, sub_838_carry_4_, sub_838_carry_5_,
         sub_838_carry_6_, sub_832_carry_2_, sub_832_carry_3_,
         sub_832_carry_4_, sub_832_carry_5_, sub_832_carry_6_,
         sub_826_carry_2_, sub_826_carry_3_, sub_826_carry_4_,
         sub_826_carry_5_, sub_826_carry_6_, sub_820_carry_2_,
         sub_820_carry_3_, sub_820_carry_4_, sub_820_carry_5_,
         sub_820_carry_6_, sub_817_carry_2_, sub_817_carry_3_,
         sub_817_carry_4_, sub_817_carry_5_, sub_817_carry_6_, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634;
  wire   [1:0] current_state;
  wire   [1:0] next_state;
  wire   [5:0] count_state_idle;
  wire   [7:0] next;
  wire   [3:1] reg_matrix_size;
  wire   [15:0] count;
  wire   [3:0] temp_i_mat_idx;
  wire   [3:0] temp_w_mat_idx;
  wire   [8:0] reg_invalid2;
  wire   [6:0] A1;
  wire   [6:0] count08;
  wire   [6:0] count18;
  wire   [6:0] count28;
  wire   [6:0] count38;
  wire   [6:0] count48;
  wire   [6:0] count58;
  wire   [6:0] count68;
  wire   [6:0] count78;
  wire   [6:0] A3;
  wire   [127:0] D1;
  wire   [15:0] D3;
  wire   [39:0] y_out_sum0;
  wire   [39:0] y_out_sum1;
  wire   [39:0] y_out_sum2;
  wire   [39:0] y_out_sum3;
  wire   [39:0] y_out_sum4;
  wire   [39:0] y_out_sum5;
  wire   [39:0] y_out_sum6;
  wire   [39:0] y_out_sum7;
  wire   [39:0] y_out_sum8;
  wire   [39:0] y_out_sum9;
  wire   [39:0] y_out_sum10;
  wire   [39:0] y_out_sum11;
  wire   [39:0] y_out_sum12;
  wire   [39:0] y_out_sum13;
  wire   [39:0] y_out_sum14;
  wire   [39:0] sum;
  wire   [5:0] length1;
  wire   [5:0] length2;
  wire   [5:0] length3;
  wire   [5:0] length4;
  wire   [5:0] length5;
  wire   [5:0] length6;
  wire   [5:0] length7;
  wire   [5:0] length8;
  wire   [5:0] length9;
  wire   [5:0] length10;
  wire   [5:0] length11;
  wire   [5:0] length12;
  wire   [5:0] length13;
  wire   [5:0] length14;
  wire   [5:0] reg_length0;
  wire   [5:0] reg_length1;
  wire   [5:0] shift;
  wire   [5:0] reg_length2;
  wire   [5:0] reg_length3;
  wire   [5:0] reg_length4;
  wire   [5:0] reg_length5;
  wire   [5:0] reg_length6;
  wire   [5:0] reg_length7;
  wire   [5:0] reg_length8;
  wire   [5:0] reg_length9;
  wire   [5:0] reg_length10;
  wire   [5:0] reg_length11;
  wire   [5:0] reg_length12;
  wire   [5:0] reg_length13;
  wire   [5:0] reg_length14;
  wire   [5:3] reg_length00;
  wire   [5:1] reg_length01;
  wire   [5:1] reg_length02;
  wire   [5:1] reg_length03;
  wire   [5:1] reg_length04;
  wire   [5:1] reg_length05;
  wire   [5:0] reg_length06;
  wire   [5:0] reg_length07;
  wire   [5:0] reg_length08;
  wire   [5:0] reg_length09;
  wire   [5:0] reg_length010;
  wire   [5:0] reg_length011;
  wire   [5:0] reg_length012;
  wire   [5:0] reg_length013;
  wire   [5:0] reg_length014;
  wire   [2:0] count1;
  wire   [2:0] count2;
  wire   [2:0] count3;
  wire   [2:0] count4;
  wire   [2:0] count5;
  wire   [2:0] count6;
  wire   [2:0] count7;
  wire   [2:0] count8;
  wire   [2:0] count9;
  wire   [2:0] count10;
  wire   [2:0] count11;
  wire   [2:0] count12;
  wire   [2:0] count13;
  wire   [2:0] count14;
  wire   [15:0] w_in0;
  wire   [15:0] w_in1;
  wire   [15:0] w_in2;
  wire   [15:0] w_in3;
  wire   [15:0] w_in4;
  wire   [15:0] w_in5;
  wire   [15:0] w_in6;
  wire   [15:0] w_in7;
  wire   [15:0] x_in0;
  wire   [15:0] x_in1;
  wire   [15:0] x_in2;
  wire   [15:0] x_in3;
  wire   [15:0] x_in4;
  wire   [15:0] x_in5;
  wire   [15:0] x_in6;
  wire   [15:0] x_in7;
  wire   [6:3] sub_841_carry;
  wire   [6:3] sub_829_carry;
  wire   [5:2] r889_carry;
  tri   [15:0] store_matrix0;
  tri   [15:0] store_matrix1;
  tri   [15:0] store_matrix2;
  tri   [15:0] store_matrix3;
  tri   [15:0] store_matrix4;
  tri   [15:0] store_matrix5;
  tri   [15:0] store_matrix6;
  tri   [15:0] store_matrix7;
  tri   [15:0] Q02;
  tri   [15:0] Q12;
  tri   [15:0] Q22;
  tri   [15:0] Q32;
  tri   [15:0] Q42;
  tri   [15:0] Q52;
  tri   [15:0] Q62;
  tri   [15:0] Q72;

  RA1SH inst_RA1SH0 ( .Q({store_matrix0, store_matrix1, store_matrix2, 
        store_matrix3, store_matrix4, store_matrix5, store_matrix6, 
        store_matrix7}), .A(A1), .D(D1), .CLK(clk), .CEN(1'b0), .OEN(1'b0), 
        .WEN(N11045) );
  RA2SH inst_RA2SH0 ( .Q(Q02), .A({n5367, n5368, n5369, n5370, n5371, n5372, 
        n5366}), .D(D3), .CLK(clk), .CEN(1'b0), .OEN(1'b0), .WEN(WEN03) );
  RA2SH inst_RA2SH1 ( .Q(Q12), .A({n5367, n5368, n5369, n5370, n5371, n5372, 
        n5366}), .D(D3), .CLK(clk), .CEN(1'b0), .OEN(1'b0), .WEN(WEN13) );
  RA2SH inst_RA2SH2 ( .Q(Q22), .A({n5367, n5368, n5369, n5370, n5371, n5372, 
        n5366}), .D(D3), .CLK(clk), .CEN(1'b0), .OEN(1'b0), .WEN(WEN23) );
  RA2SH inst_RA2SH3 ( .Q(Q32), .A({n5367, n5368, n5369, n5370, n5371, n5372, 
        n5366}), .D(D3), .CLK(clk), .CEN(1'b0), .OEN(1'b0), .WEN(WEN33) );
  RA2SH inst_RA2SH4 ( .Q(Q42), .A({n5367, n5368, n5369, n5370, n5371, n5372, 
        n5366}), .D(D3), .CLK(clk), .CEN(1'b0), .OEN(1'b0), .WEN(WEN43) );
  RA2SH inst_RA2SH5 ( .Q(Q52), .A({n5367, n5368, n5369, n5370, n5371, n5372, 
        n5366}), .D(D3), .CLK(clk), .CEN(1'b0), .OEN(1'b0), .WEN(WEN53) );
  RA2SH inst_RA2SH6 ( .Q(Q62), .A({n5367, n5368, n5369, n5370, n5371, n5372, 
        n5366}), .D(D3), .CLK(clk), .CEN(1'b0), .OEN(1'b0), .WEN(WEN63) );
  RA2SH inst_RA2SH7 ( .Q(Q72), .A({n5367, n5368, n5369, n5370, n5371, n5372, 
        n5366}), .D(D3), .CLK(clk), .CEN(1'b0), .OEN(1'b0), .WEN(WEN73) );
  DFFHQX4 w_in7_reg_9_ ( .D(n7136), .CK(clk), .Q(w_in7[9]) );
  DFFHQX4 w_in7_reg_7_ ( .D(n7138), .CK(clk), .Q(w_in7[7]) );
  DFFHQX4 w_in3_reg_9_ ( .D(n3009), .CK(clk), .Q(w_in3[9]) );
  DFFHQX4 w_in3_reg_7_ ( .D(n3011), .CK(clk), .Q(w_in3[7]) );
  DFFHQX4 w_in7_reg_5_ ( .D(n7140), .CK(clk), .Q(w_in7[5]) );
  DFFHQX4 w_in3_reg_5_ ( .D(n3013), .CK(clk), .Q(w_in3[5]) );
  DFFHQX4 w_in4_reg_3_ ( .D(n3111), .CK(clk), .Q(w_in4[3]) );
  DFFHQX4 w_in4_reg_1_ ( .D(n3113), .CK(clk), .Q(w_in4[1]) );
  DFFHQX4 w_in7_reg_3_ ( .D(n7142), .CK(clk), .Q(w_in7[3]) );
  DFFHQX4 w_in3_reg_3_ ( .D(n3015), .CK(clk), .Q(w_in3[3]) );
  DFFHQX4 w_in5_reg_5_ ( .D(n3093), .CK(clk), .Q(w_in5[5]) );
  DFFHQX4 w_in5_reg_3_ ( .D(n3095), .CK(clk), .Q(w_in5[3]) );
  DFFHQX4 w_in5_reg_1_ ( .D(n3097), .CK(clk), .Q(w_in5[1]) );
  DFFHQX4 w_in2_reg_13_ ( .D(n3069), .CK(clk), .Q(w_in2[13]) );
  DFFHQX4 w_in6_reg_11_ ( .D(n7148), .CK(clk), .Q(w_in6[11]) );
  DFFHQX4 w_in2_reg_11_ ( .D(n3071), .CK(clk), .Q(w_in2[11]) );
  DFFHQX4 w_in2_reg_9_ ( .D(n3073), .CK(clk), .Q(w_in2[9]) );
  DFFHQX4 w_in2_reg_7_ ( .D(n3075), .CK(clk), .Q(w_in2[7]) );
  DFFHQX4 w_in6_reg_5_ ( .D(n7154), .CK(clk), .Q(w_in6[5]) );
  DFFHQX4 w_in2_reg_5_ ( .D(n3077), .CK(clk), .Q(w_in2[5]) );
  DFFHQX4 w_in7_reg_1_ ( .D(n7156), .CK(clk), .Q(w_in7[1]) );
  DFFHQX4 w_in1_reg_1_ ( .D(n3033), .CK(clk), .Q(w_in1[1]) );
  DFFHQX4 w_in3_reg_1_ ( .D(n3017), .CK(clk), .Q(w_in3[1]) );
  DFFHQX4 w_in6_reg_3_ ( .D(n7157), .CK(clk), .Q(w_in6[3]) );
  DFFHQX4 w_in2_reg_3_ ( .D(n3079), .CK(clk), .Q(w_in2[3]) );
  DFFHQX4 w_in6_reg_1_ ( .D(n7159), .CK(clk), .Q(w_in6[1]) );
  DFFHQX4 w_in2_reg_1_ ( .D(n3081), .CK(clk), .Q(w_in2[1]) );
  DFFHQX4 w_in3_reg_13_ ( .D(n3005), .CK(clk), .Q(w_in3[13]) );
  DFFHQX4 w_in0_reg_13_ ( .D(n3037), .CK(clk), .Q(w_in0[13]) );
  DFFHQX4 w_in0_reg_11_ ( .D(n3039), .CK(clk), .Q(w_in0[11]) );
  DFFHQX4 w_in0_reg_9_ ( .D(n3041), .CK(clk), .Q(w_in0[9]) );
  DFFHQX4 w_in3_reg_11_ ( .D(n3007), .CK(clk), .Q(w_in3[11]) );
  DFFHQX4 w_in0_reg_7_ ( .D(n3043), .CK(clk), .Q(w_in0[7]) );
  DFFHQX4 w_in0_reg_5_ ( .D(n3045), .CK(clk), .Q(w_in0[5]) );
  DFFHQX4 w_in0_reg_3_ ( .D(n3047), .CK(clk), .Q(w_in0[3]) );
  DFFHQX4 w_in0_reg_1_ ( .D(n3049), .CK(clk), .Q(w_in0[1]) );
  DFFHQX4 w_in1_reg_13_ ( .D(n3021), .CK(clk), .Q(w_in1[13]) );
  DFFHQX4 w_in1_reg_11_ ( .D(n3023), .CK(clk), .Q(w_in1[11]) );
  DFFHQX4 w_in1_reg_9_ ( .D(n3025), .CK(clk), .Q(w_in1[9]) );
  DFFHQX4 w_in1_reg_7_ ( .D(n3027), .CK(clk), .Q(w_in1[7]) );
  compare_0 inst_compare1 ( .clk(clk), .rst(1'b0), .sum(y_out_sum1), .length(
        length1) );
  compare_13 inst_compare2 ( .clk(clk), .rst(1'b0), .sum(y_out_sum2), .length(
        length2) );
  compare_12 inst_compare3 ( .clk(clk), .rst(1'b0), .sum(y_out_sum3), .length(
        length3) );
  compare_11 inst_compare4 ( .clk(clk), .rst(1'b0), .sum(y_out_sum4), .length(
        length4) );
  compare_10 inst_compare5 ( .clk(clk), .rst(1'b0), .sum(y_out_sum5), .length(
        length5) );
  compare_9 inst_compare6 ( .clk(clk), .rst(1'b0), .sum(y_out_sum6), .length(
        length6) );
  compare_8 inst_compare7 ( .clk(clk), .rst(1'b0), .sum(y_out_sum7), .length(
        length7) );
  compare_7 inst_compare8 ( .clk(clk), .rst(1'b0), .sum(y_out_sum8), .length(
        length8) );
  compare_6 inst_compare9 ( .clk(clk), .rst(1'b0), .sum(y_out_sum9), .length(
        length9) );
  compare_5 inst_compare10 ( .clk(clk), .rst(1'b0), .sum(y_out_sum10), 
        .length(length10) );
  compare_4 inst_compare11 ( .clk(clk), .rst(1'b0), .sum(y_out_sum11), 
        .length(length11) );
  compare_3 inst_compare12 ( .clk(clk), .rst(1'b0), .sum(y_out_sum12), 
        .length(length12) );
  compare_2 inst_compare13 ( .clk(clk), .rst(1'b0), .sum(y_out_sum13), 
        .length(length13) );
  compare_1 inst_compare14 ( .clk(clk), .rst(1'b0), .sum(y_out_sum14), 
        .length(length14) );
  PE inst_PE ( .clk(clk), .rst(1'b0), .x_in0(x_in0), .x_in1(x_in1), .x_in2(
        x_in2), .x_in3(x_in3), .x_in4(x_in4), .x_in5(x_in5), .x_in6(x_in6), 
        .x_in7(x_in7), .w_in0(w_in0), .w_in1(w_in1), .w_in2(w_in2), .w_in3(
        w_in3), .w_in4(w_in4), .w_in5(w_in5), .w_in6(w_in6), .w_in7(w_in7), 
        .y_out(sum) );
  MMSA_DW01_inc_0_DW01_inc_14 add_738 ( .A(count78), .SUM({N4969, N4968, N4967, 
        N4966, N4965, N4964, N4963}) );
  MMSA_DW01_inc_1_DW01_inc_15 add_724 ( .A(count68), .SUM({N4952, N4951, N4950, 
        N4949, N4948, N4947, N4946}) );
  MMSA_DW01_inc_2_DW01_inc_16 add_710 ( .A(count58), .SUM({N4935, N4934, N4933, 
        N4932, N4931, N4930, N4929}) );
  MMSA_DW01_inc_3_DW01_inc_17 add_696 ( .A(count48), .SUM({N4918, N4917, N4916, 
        N4915, N4914, N4913, N4912}) );
  MMSA_DW01_inc_4_DW01_inc_18 add_682 ( .A(count38), .SUM({N4901, N4900, N4899, 
        N4898, N4897, N4896, N4895}) );
  MMSA_DW01_inc_5_DW01_inc_19 add_668 ( .A(count28), .SUM({N4884, N4883, N4882, 
        N4881, N4880, N4879, N4878}) );
  MMSA_DW01_inc_6_DW01_inc_20 add_654 ( .A(count18), .SUM({N4867, N4866, N4865, 
        N4864, N4863, N4862, N4861}) );
  MMSA_DW01_inc_7_DW01_inc_21 add_640 ( .A(count08), .SUM({N4850, N4849, N4848, 
        N4847, N4846, N4845, N4844}) );
  MMSA_DW01_inc_8_DW01_inc_22 add_248 ( .A({count[15:13], n5377, n5378, N5118, 
        n5568, N5061, n5571, N5059, n5379, n5380, count[3:0]}), .SUM({N4599, 
        N4598, N4597, N4596, N4595, N4594, N4593, N4592, N4591, N4590, N4589, 
        N4588, N4587, N4586, N4585, N4584}) );
  MMSA_DW01_inc_9_DW01_inc_23 r964 ( .A(next), .SUM({N8524, N8523, N8522, 
        N8521, N8520, N8519, N8518, N8517}) );
  MMSA_DW01_inc_10_DW01_inc_24 r892 ( .A({reg_invalid2[8:6], n5373, 
        reg_invalid2[4], n5374, n5375, n5376, reg_invalid2[0]}), .SUM({N4702, 
        N4701, N4700, N4699, N4698, N4697, N4696, N4695, N4694}) );
  MMSA_DW01_add_30 add_1067 ( .A(y_out_sum14), .B({sum[39], n5556, n5560, 
        n4843, n5565, n5553, n5551, n5347, n5547, n5545, n5543, n5541, n5539, 
        n5536, n4846, n5531, n5529, n5527, n5525, n5523, n4983, n5518, n4978, 
        n5514, n4844, n5509, n5507, n5505, n5502, n5499, n5497, n5495, n5492, 
        n5489, n4967, n5484, n5481, n5479, n5476, n5474}), .CI(1'b0), .SUM({
        N6497, N6496, N6495, N6494, N6493, N6492, N6491, N6490, N6489, N6488, 
        N6487, N6486, N6485, N6484, N6483, N6482, N6481, N6480, N6479, N6478, 
        N6477, N6476, N6475, N6474, N6473, N6472, N6471, N6470, N6469, N6468, 
        N6467, N6466, N6465, N6464, N6463, N6462, N6461, N6460, N6459, N6458})
         );
  MMSA_DW01_add_31 add_1064 ( .A(y_out_sum13), .B({sum[39], n5556, n5560, 
        n4843, n5565, sum[34], n5551, n5347, n5547, n5545, n5543, n4972, n4975, 
        n5536, n4846, n5531, n5529, n5527, n5525, n5523, n4983, n4986, n4978, 
        n5514, n5511, n5509, n5507, n5505, n5502, n5499, n5497, n5495, n5492, 
        n4971, n4967, n5484, n5481, n5479, n5476, sum[0]}), .CI(1'b0), .SUM({
        N6456, N6455, N6454, N6453, N6452, N6451, N6450, N6449, N6448, N6447, 
        N6446, N6445, N6444, N6443, N6442, N6441, N6440, N6439, N6438, N6437, 
        N6436, N6435, N6434, N6433, N6432, N6431, N6430, N6429, N6428, N6427, 
        N6426, N6425, N6424, N6423, N6422, N6421, N6420, N6419, N6418, N6417})
         );
  MMSA_DW01_add_32 add_1061 ( .A(y_out_sum12), .B({sum[39], n5555, n5560, 
        n4843, n5565, sum[34], n5551, n5347, n5547, n4982, n5543, n5541, n4975, 
        n5536, sum[25], n5531, n4976, n5527, sum[21], n5523, n5521, n4985, 
        n5516, n5514, n5511, n5509, n4969, n5505, n5502, n5499, n5497, n5495, 
        n5492, n5489, n5487, n5484, n5481, sum[2], n5476, sum[0]}), .CI(1'b0), 
        .SUM({N6415, N6414, N6413, N6412, N6411, N6410, N6409, N6408, N6407, 
        N6406, N6405, N6404, N6403, N6402, N6401, N6400, N6399, N6398, N6397, 
        N6396, N6395, N6394, N6393, N6392, N6391, N6390, N6389, N6388, N6387, 
        N6386, N6385, N6384, N6383, N6382, N6381, N6380, N6379, N6378, N6377, 
        N6376}) );
  MMSA_DW01_add_33 add_1058 ( .A(y_out_sum11), .B({sum[39], n5555, n5559, 
        n4843, n4843, n5553, n5551, n5549, n5547, n4974, n5543, n5541, n5539, 
        n5535, n4846, n5531, n4977, n5527, n5525, n5523, n5521, n4985, n4978, 
        n5513, n4844, n5509, n4969, n5504, n5502, n5499, n5497, n5495, n5492, 
        n4971, n5487, n5484, n5481, n5479, n5476, n5474}), .CI(1'b0), .SUM({
        N6374, N6373, N6372, N6371, N6370, N6369, N6368, N6367, N6366, N6365, 
        N6364, N6363, N6362, N6361, N6360, N6359, N6358, N6357, N6356, N6355, 
        N6354, N6353, N6352, N6351, N6350, N6349, N6348, N6347, N6346, N6345, 
        N6344, N6343, N6342, N6341, N6340, N6339, N6338, N6337, N6336, N6335})
         );
  MMSA_DW01_add_34 add_1055 ( .A(y_out_sum10), .B({sum[39], n5555, n4984, 
        n4843, n4843, n5553, n5551, n5549, n5547, n4982, n5543, n4972, n5538, 
        n5535, n4846, n5531, n4976, n5527, n5525, n5523, n5521, n4985, n5516, 
        n5513, n5511, n5509, n5507, n5504, n5502, n5499, n5497, n5495, n5492, 
        n5489, n5487, n5484, n5481, n5479, n5476, n5474}), .CI(1'b0), .SUM({
        N6333, N6332, N6331, N6330, N6329, N6328, N6327, N6326, N6325, N6324, 
        N6323, N6322, N6321, N6320, N6319, N6318, N6317, N6316, N6315, N6314, 
        N6313, N6312, N6311, N6310, N6309, N6308, N6307, N6306, N6305, N6304, 
        N6303, N6302, N6301, N6300, N6299, N6298, N6297, N6296, N6295, N6294})
         );
  MMSA_DW01_add_35 add_1052 ( .A(y_out_sum9), .B({sum[39], n5555, n4984, n4843, 
        n4841, n5553, n5551, n5347, n5547, n4974, n5543, n4972, n5538, n5535, 
        n4846, n5531, sum[23], n5527, n5525, n5523, n4983, n4986, sum[17], 
        n5513, n5511, n5509, n4968, n5504, n5502, n5499, n5497, n5495, n5492, 
        n5490, n4967, n5484, n5481, n5479, n5476, n5474}), .CI(1'b0), .SUM({
        N6292, N6291, N6290, N6289, N6288, N6287, N6286, N6285, N6284, N6283, 
        N6282, N6281, N6280, N6279, N6278, N6277, N6276, N6275, N6274, N6273, 
        N6272, N6271, N6270, N6269, N6268, N6267, N6266, N6265, N6264, N6263, 
        N6262, N6261, N6260, N6259, N6258, N6257, N6256, N6255, N6254, N6253})
         );
  MMSA_DW01_add_36 add_1049 ( .A(y_out_sum8), .B({sum[39], n5555, n4984, n4843, 
        n4843, n5553, n5551, n5549, n5547, n4974, n5543, n5541, sum[27], n5535, 
        n4846, n5531, n5529, n5527, n5525, n5523, n4983, n4985, n5516, n5513, 
        n4844, n5509, n4968, n5504, n5502, n5499, n5497, n5495, n5492, n5489, 
        n4967, n5484, n5481, n5479, n5476, n5474}), .CI(1'b0), .SUM({N6251, 
        N6250, N6249, N6248, N6247, N6246, N6245, N6244, N6243, N6242, N6241, 
        N6240, N6239, N6238, N6237, N6236, N6235, N6234, N6233, N6232, N6231, 
        N6230, N6229, N6228, N6227, N6226, N6225, N6224, N6223, N6222, N6221, 
        N6220, N6219, N6218, N6217, N6216, N6215, N6214, N6213, N6212}) );
  MMSA_DW01_add_37 add_1046 ( .A(y_out_sum7), .B({sum[39], n5555, n4984, n4843, 
        n4843, n5553, n5551, n5347, n5547, n4982, n5543, n4972, n5538, n5535, 
        n4846, n5531, n4977, n5527, n5525, n5523, n4983, n4986, n4978, sum[16], 
        n5511, n5509, n4969, n5504, n5502, n5499, n5497, n5495, n5492, n5490, 
        n4967, n5484, n5481, n5479, n5476, n5474}), .CI(1'b0), .SUM({N6210, 
        N6209, N6208, N6207, N6206, N6205, N6204, N6203, N6202, N6201, N6200, 
        N6199, N6198, N6197, N6196, N6195, N6194, N6193, N6192, N6191, N6190, 
        N6189, N6188, N6187, N6186, N6185, N6184, N6183, N6182, N6181, N6180, 
        N6179, N6178, N6177, N6176, N6175, N6174, N6173, N6172, N6171}) );
  MMSA_DW01_add_38 r924 ( .A(y_out_sum6), .B({sum[39], n5555, n5559, n4843, 
        n5565, n4842, n5551, n5347, n5547, n5545, n5543, n5541, sum[27], n5535, 
        n4846, n5531, n5529, n5527, n5525, n5523, n5520, n4985, n5516, sum[16], 
        n5511, n5509, n5507, n5504, n5502, n5499, n5497, n5495, n5492, n5490, 
        n5487, n5484, n5481, n5479, n5476, n5474}), .CI(1'b0), .SUM({N5845, 
        N5844, N5843, N5842, N5841, N5840, N5839, N5838, N5837, N5836, N5835, 
        N5834, N5833, N5832, N5831, N5830, N5829, N5828, N5827, N5826, N5825, 
        N5824, N5823, N5822, N5821, N5820, N5819, N5818, N5817, N5816, N5815, 
        N5814, N5813, N5812, N5811, N5810, N5809, N5808, N5807, N5806}) );
  MMSA_DW01_add_39 r923 ( .A(y_out_sum5), .B({sum[39], n5555, n5559, n4843, 
        n4841, n4842, n5551, n5347, n5547, n5545, n5543, n5541, sum[27], n5535, 
        n4846, n5531, n4976, n5527, n5525, n5523, n5521, n5518, n4978, n5513, 
        n5511, n5509, n4968, n5504, n5502, n5499, n5497, n5495, n5492, n5489, 
        n4967, n5484, n5481, n5479, n5476, n5474}), .CI(1'b0), .SUM({N5804, 
        N5803, N5802, N5801, N5800, N5799, N5798, N5797, N5796, N5795, N5794, 
        N5793, N5792, N5791, N5790, N5789, N5788, N5787, N5786, N5785, N5784, 
        N5783, N5782, N5781, N5780, N5779, N5778, N5777, N5776, N5775, N5774, 
        N5773, N5772, N5771, N5770, N5769, N5768, N5767, N5766, N5765}) );
  MMSA_DW01_add_40 r922 ( .A(y_out_sum4), .B({sum[39], n5555, n5559, n4842, 
        n4841, n4842, n5551, n5549, n5547, n5545, n5543, n4972, n5538, n5535, 
        n4845, n5531, n5529, n5527, n5525, n5523, n5520, n5518, n5516, sum[16], 
        n5511, n5509, n5507, n5504, n5502, n5499, n5497, n5495, n5492, n5490, 
        n5487, n5484, n5481, n5479, n5476, n5474}), .CI(1'b0), .SUM({N5763, 
        N5762, N5761, N5760, N5759, N5758, N5757, N5756, N5755, N5754, N5753, 
        N5752, N5751, N5750, N5749, N5748, N5747, N5746, N5745, N5744, N5743, 
        N5742, N5741, N5740, N5739, N5738, N5737, N5736, N5735, N5734, N5733, 
        N5732, N5731, N5730, N5729, N5728, N5727, N5726, N5725, N5724}) );
  MMSA_DW01_add_41 r921 ( .A(y_out_sum3), .B({sum[39], n5555, n5559, n4843, 
        n4841, n4842, n5551, n5347, n5547, n5545, n5543, n5541, n5538, n5535, 
        n4846, n5531, n5529, n5527, n5525, n5523, n4983, n4985, n4978, sum[16], 
        n5511, n5509, n4969, n5504, n5502, n5500, sum[9], n5495, n5493, n4971, 
        n5487, n5485, n5482, n5479, n5477, n5474}), .CI(1'b0), .SUM({N5722, 
        N5721, N5720, N5719, N5718, N5717, N5716, N5715, N5714, N5713, N5712, 
        N5711, N5710, N5709, N5708, N5707, N5706, N5705, N5704, N5703, N5702, 
        N5701, N5700, N5699, N5698, N5697, N5696, N5695, N5694, N5693, N5692, 
        N5691, N5690, N5689, N5688, N5687, N5686, N5685, N5684, N5683}) );
  MMSA_DW01_add_42 r920 ( .A(y_out_sum2), .B({sum[39], n5555, n5559, n4843, 
        n4841, n4842, n5551, n5347, n5547, n5545, n5543, n4972, sum[27], n5535, 
        n4846, n5531, n4976, n5527, n5525, n5523, n5520, n5518, n5516, sum[16], 
        n5511, n5509, n4968, n5504, n5502, n5500, sum[9], n5495, n5493, n5489, 
        n4967, n5485, n5482, n5479, n5477, n5474}), .CI(1'b0), .SUM({N5541, 
        N5540, N5539, N5538, N5537, N5536, N5535, N5534, N5533, N5532, N5531, 
        N5530, N5529, N5528, N5527, N5526, N5525, N5524, N5523, N5522, N5521, 
        N5520, N5519, N5518, N5517, N5516, N5515, N5514, N5513, N5512, N5511, 
        N5510, N5509, N5508, N5507, N5506, N5505, N5504, N5503, N5502}) );
  MMSA_DW01_add_43 r919 ( .A(y_out_sum1), .B({sum[39], n5555, n5559, n4843, 
        n4840, n4842, n5551, n5347, n5547, n5545, n5543, n4972, sum[27], n5535, 
        n4846, n5531, n4977, n5527, n5525, n5523, n5520, n4985, n4978, sum[16], 
        n4844, n5509, n4968, n5504, n5502, n5500, n5497, n5495, n5493, n4971, 
        n5487, n5485, n5482, n5479, n5477, n5474}), .CI(1'b0), .SUM({N5500, 
        N5499, N5498, N5497, N5496, N5495, N5494, N5493, N5492, N5491, N5490, 
        N5489, N5488, N5487, N5486, N5485, N5484, N5483, N5482, N5481, N5480, 
        N5479, N5478, N5477, N5476, N5475, N5474, N5473, N5472, N5471, N5470, 
        N5469, N5468, N5467, N5466, N5465, N5464, N5463, N5462, N5461}) );
  MMSA_DW01_add_44 r918 ( .A(y_out_sum0), .B({sum[39], n5555, n5559, n4843, 
        n4841, n5553, n5551, n5347, n5547, n4973, n5543, n5541, n4975, n5535, 
        n4846, n5531, n4977, n5527, n5525, n5523, n5521, n4986, n5516, n5513, 
        n5511, n5509, n4968, n5504, n5502, n5499, n5497, n5495, n5492, n4971, 
        n4967, n5484, n5481, n5479, n5476, n5474}), .CI(1'b0), .SUM({N5459, 
        N5458, N5457, N5456, N5455, N5454, N5453, N5452, N5451, N5450, N5449, 
        N5448, N5447, N5446, N5445, N5444, N5443, N5442, N5441, N5440, N5439, 
        N5438, N5437, N5436, N5435, N5434, N5433, N5432, N5431, N5430, N5429, 
        N5428, N5427, N5426, N5425, N5424, N5423, N5422, N5421, N5420}) );
  DFFX4 w_in6_reg_9_ ( .D(n7150), .CK(clk), .Q(w_in6[9]), .QN(n5600) );
  DFFX4 w_in4_reg_7_ ( .D(n3107), .CK(clk), .Q(w_in4[7]), .QN(n5630) );
  DFFX4 w_in4_reg_5_ ( .D(n3109), .CK(clk), .Q(w_in4[5]), .QN(n5628) );
  DFFRXL y_out_sum9_reg_39_ ( .D(n3506), .CK(clk), .RN(rst_n), .Q(
        y_out_sum9[39]), .QN(n6662) );
  DFFRHQX1 D1_reg_0_ ( .D(N5258), .CK(clk), .RN(rst_n), .Q(D1[0]) );
  DFFRHQX1 D1_reg_1_ ( .D(N5259), .CK(clk), .RN(rst_n), .Q(D1[1]) );
  DFFRHQX1 D1_reg_2_ ( .D(N5260), .CK(clk), .RN(rst_n), .Q(D1[2]) );
  DFFRHQX1 D1_reg_3_ ( .D(N5261), .CK(clk), .RN(rst_n), .Q(D1[3]) );
  DFFRHQX1 D1_reg_4_ ( .D(N5262), .CK(clk), .RN(rst_n), .Q(D1[4]) );
  DFFRHQX1 D1_reg_5_ ( .D(N5263), .CK(clk), .RN(rst_n), .Q(D1[5]) );
  DFFRHQX1 D1_reg_6_ ( .D(N5264), .CK(clk), .RN(rst_n), .Q(D1[6]) );
  DFFRHQX1 D1_reg_7_ ( .D(N5265), .CK(clk), .RN(rst_n), .Q(D1[7]) );
  DFFRHQX1 D1_reg_8_ ( .D(N5266), .CK(clk), .RN(rst_n), .Q(D1[8]) );
  DFFRHQX1 D1_reg_9_ ( .D(N5267), .CK(clk), .RN(rst_n), .Q(D1[9]) );
  DFFRHQX1 D1_reg_10_ ( .D(N5268), .CK(clk), .RN(rst_n), .Q(D1[10]) );
  DFFRHQX1 D1_reg_11_ ( .D(N5269), .CK(clk), .RN(rst_n), .Q(D1[11]) );
  DFFRHQX1 D1_reg_12_ ( .D(N5270), .CK(clk), .RN(rst_n), .Q(D1[12]) );
  DFFRHQX1 D1_reg_13_ ( .D(N5271), .CK(clk), .RN(rst_n), .Q(D1[13]) );
  DFFRHQX1 D1_reg_14_ ( .D(N5272), .CK(clk), .RN(rst_n), .Q(D1[14]) );
  DFFRHQX1 D1_reg_15_ ( .D(N5273), .CK(clk), .RN(rst_n), .Q(D1[15]) );
  DFFRHQX1 D1_reg_16_ ( .D(N5274), .CK(clk), .RN(rst_n), .Q(D1[16]) );
  DFFRHQX1 D1_reg_17_ ( .D(N5275), .CK(clk), .RN(rst_n), .Q(D1[17]) );
  DFFRHQX1 D1_reg_18_ ( .D(N5276), .CK(clk), .RN(rst_n), .Q(D1[18]) );
  DFFRHQX1 D1_reg_19_ ( .D(N5277), .CK(clk), .RN(rst_n), .Q(D1[19]) );
  DFFRHQX1 D1_reg_20_ ( .D(N5278), .CK(clk), .RN(rst_n), .Q(D1[20]) );
  DFFRHQX1 D1_reg_21_ ( .D(N5279), .CK(clk), .RN(rst_n), .Q(D1[21]) );
  DFFRHQX1 D1_reg_22_ ( .D(N5280), .CK(clk), .RN(rst_n), .Q(D1[22]) );
  DFFRHQX1 D1_reg_23_ ( .D(N5281), .CK(clk), .RN(rst_n), .Q(D1[23]) );
  DFFRHQX1 D1_reg_24_ ( .D(N5282), .CK(clk), .RN(rst_n), .Q(D1[24]) );
  DFFRHQX1 D1_reg_25_ ( .D(N5283), .CK(clk), .RN(rst_n), .Q(D1[25]) );
  DFFRHQX1 D1_reg_26_ ( .D(N5284), .CK(clk), .RN(rst_n), .Q(D1[26]) );
  DFFRHQX1 D1_reg_27_ ( .D(N5285), .CK(clk), .RN(rst_n), .Q(D1[27]) );
  DFFRHQX1 D1_reg_28_ ( .D(N5286), .CK(clk), .RN(rst_n), .Q(D1[28]) );
  DFFRHQX1 D1_reg_29_ ( .D(N5287), .CK(clk), .RN(rst_n), .Q(D1[29]) );
  DFFRHQX1 D1_reg_30_ ( .D(N5288), .CK(clk), .RN(rst_n), .Q(D1[30]) );
  DFFRHQX1 D1_reg_31_ ( .D(N5289), .CK(clk), .RN(rst_n), .Q(D1[31]) );
  DFFRHQX1 D1_reg_32_ ( .D(N5290), .CK(clk), .RN(rst_n), .Q(D1[32]) );
  DFFRHQX1 D1_reg_33_ ( .D(N5291), .CK(clk), .RN(rst_n), .Q(D1[33]) );
  DFFRHQX1 D1_reg_34_ ( .D(N5292), .CK(clk), .RN(rst_n), .Q(D1[34]) );
  DFFRHQX1 D1_reg_35_ ( .D(N5293), .CK(clk), .RN(rst_n), .Q(D1[35]) );
  DFFRHQX1 D1_reg_36_ ( .D(N5294), .CK(clk), .RN(rst_n), .Q(D1[36]) );
  DFFRHQX1 D1_reg_37_ ( .D(N5295), .CK(clk), .RN(rst_n), .Q(D1[37]) );
  DFFRHQX1 D1_reg_38_ ( .D(N5296), .CK(clk), .RN(rst_n), .Q(D1[38]) );
  DFFRHQX1 D1_reg_39_ ( .D(N5297), .CK(clk), .RN(rst_n), .Q(D1[39]) );
  DFFRHQX1 D1_reg_40_ ( .D(N5298), .CK(clk), .RN(rst_n), .Q(D1[40]) );
  DFFRHQX1 D1_reg_41_ ( .D(N5299), .CK(clk), .RN(rst_n), .Q(D1[41]) );
  DFFRHQX1 D1_reg_42_ ( .D(N5300), .CK(clk), .RN(rst_n), .Q(D1[42]) );
  DFFRHQX1 D1_reg_43_ ( .D(N5301), .CK(clk), .RN(rst_n), .Q(D1[43]) );
  DFFRHQX1 D1_reg_44_ ( .D(N5302), .CK(clk), .RN(rst_n), .Q(D1[44]) );
  DFFRHQX1 D1_reg_45_ ( .D(N5303), .CK(clk), .RN(rst_n), .Q(D1[45]) );
  DFFRHQX1 D1_reg_46_ ( .D(N5304), .CK(clk), .RN(rst_n), .Q(D1[46]) );
  DFFRHQX1 D1_reg_47_ ( .D(N5305), .CK(clk), .RN(rst_n), .Q(D1[47]) );
  DFFRHQX1 D1_reg_48_ ( .D(N5306), .CK(clk), .RN(rst_n), .Q(D1[48]) );
  DFFRHQX1 D1_reg_49_ ( .D(N5307), .CK(clk), .RN(rst_n), .Q(D1[49]) );
  DFFRHQX1 D1_reg_50_ ( .D(N5308), .CK(clk), .RN(rst_n), .Q(D1[50]) );
  DFFRHQX1 D1_reg_51_ ( .D(N5309), .CK(clk), .RN(rst_n), .Q(D1[51]) );
  DFFRHQX1 D1_reg_52_ ( .D(N5310), .CK(clk), .RN(rst_n), .Q(D1[52]) );
  DFFRHQX1 D1_reg_53_ ( .D(N5311), .CK(clk), .RN(rst_n), .Q(D1[53]) );
  DFFRHQX1 D1_reg_54_ ( .D(N5312), .CK(clk), .RN(rst_n), .Q(D1[54]) );
  DFFRHQX1 D1_reg_55_ ( .D(N5313), .CK(clk), .RN(rst_n), .Q(D1[55]) );
  DFFRHQX1 D1_reg_56_ ( .D(N5314), .CK(clk), .RN(rst_n), .Q(D1[56]) );
  DFFRHQX1 D1_reg_57_ ( .D(N5315), .CK(clk), .RN(rst_n), .Q(D1[57]) );
  DFFRHQX1 D1_reg_58_ ( .D(N5316), .CK(clk), .RN(rst_n), .Q(D1[58]) );
  DFFRHQX1 D1_reg_59_ ( .D(N5317), .CK(clk), .RN(rst_n), .Q(D1[59]) );
  DFFRHQX1 D1_reg_60_ ( .D(N5318), .CK(clk), .RN(rst_n), .Q(D1[60]) );
  DFFRHQX1 D1_reg_61_ ( .D(N5319), .CK(clk), .RN(rst_n), .Q(D1[61]) );
  DFFRHQX1 D1_reg_62_ ( .D(N5320), .CK(clk), .RN(rst_n), .Q(D1[62]) );
  DFFRHQX1 D1_reg_63_ ( .D(N5321), .CK(clk), .RN(rst_n), .Q(D1[63]) );
  DFFRHQX1 D1_reg_64_ ( .D(N5322), .CK(clk), .RN(rst_n), .Q(D1[64]) );
  DFFRHQX1 D1_reg_65_ ( .D(N5323), .CK(clk), .RN(rst_n), .Q(D1[65]) );
  DFFRHQX1 D1_reg_66_ ( .D(N5324), .CK(clk), .RN(rst_n), .Q(D1[66]) );
  DFFRHQX1 D1_reg_67_ ( .D(N5325), .CK(clk), .RN(rst_n), .Q(D1[67]) );
  DFFRHQX1 D1_reg_68_ ( .D(N5326), .CK(clk), .RN(rst_n), .Q(D1[68]) );
  DFFRHQX1 D1_reg_69_ ( .D(N5327), .CK(clk), .RN(rst_n), .Q(D1[69]) );
  DFFRHQX1 D1_reg_70_ ( .D(N5328), .CK(clk), .RN(rst_n), .Q(D1[70]) );
  DFFRHQX1 D1_reg_71_ ( .D(N5329), .CK(clk), .RN(rst_n), .Q(D1[71]) );
  DFFRHQX1 D1_reg_72_ ( .D(N5330), .CK(clk), .RN(rst_n), .Q(D1[72]) );
  DFFRHQX1 D1_reg_73_ ( .D(N5331), .CK(clk), .RN(rst_n), .Q(D1[73]) );
  DFFRHQX1 D1_reg_74_ ( .D(N5332), .CK(clk), .RN(rst_n), .Q(D1[74]) );
  DFFRHQX1 D1_reg_75_ ( .D(N5333), .CK(clk), .RN(rst_n), .Q(D1[75]) );
  DFFRHQX1 D1_reg_76_ ( .D(N5334), .CK(clk), .RN(rst_n), .Q(D1[76]) );
  DFFRHQX1 D1_reg_77_ ( .D(N5335), .CK(clk), .RN(rst_n), .Q(D1[77]) );
  DFFRHQX1 D1_reg_78_ ( .D(N5336), .CK(clk), .RN(rst_n), .Q(D1[78]) );
  DFFRHQX1 D1_reg_79_ ( .D(N5337), .CK(clk), .RN(rst_n), .Q(D1[79]) );
  DFFRHQX1 D1_reg_80_ ( .D(N5338), .CK(clk), .RN(rst_n), .Q(D1[80]) );
  DFFRHQX1 D1_reg_81_ ( .D(N5339), .CK(clk), .RN(rst_n), .Q(D1[81]) );
  DFFRHQX1 D1_reg_82_ ( .D(N5340), .CK(clk), .RN(rst_n), .Q(D1[82]) );
  DFFRHQX1 D1_reg_83_ ( .D(N5341), .CK(clk), .RN(rst_n), .Q(D1[83]) );
  DFFRHQX1 D1_reg_84_ ( .D(N5342), .CK(clk), .RN(rst_n), .Q(D1[84]) );
  DFFRHQX1 D1_reg_85_ ( .D(N5343), .CK(clk), .RN(rst_n), .Q(D1[85]) );
  DFFRHQX1 D1_reg_86_ ( .D(N5344), .CK(clk), .RN(rst_n), .Q(D1[86]) );
  DFFRHQX1 D1_reg_87_ ( .D(N5345), .CK(clk), .RN(rst_n), .Q(D1[87]) );
  DFFRHQX1 D1_reg_88_ ( .D(N5346), .CK(clk), .RN(rst_n), .Q(D1[88]) );
  DFFRHQX1 D1_reg_89_ ( .D(N5347), .CK(clk), .RN(rst_n), .Q(D1[89]) );
  DFFRHQX1 D1_reg_90_ ( .D(N5348), .CK(clk), .RN(rst_n), .Q(D1[90]) );
  DFFRHQX1 D1_reg_91_ ( .D(N5349), .CK(clk), .RN(rst_n), .Q(D1[91]) );
  DFFRHQX1 D1_reg_92_ ( .D(N5350), .CK(clk), .RN(rst_n), .Q(D1[92]) );
  DFFRHQX1 D1_reg_93_ ( .D(N5351), .CK(clk), .RN(rst_n), .Q(D1[93]) );
  DFFRHQX1 D1_reg_94_ ( .D(N5352), .CK(clk), .RN(rst_n), .Q(D1[94]) );
  DFFRHQX1 D1_reg_95_ ( .D(N5353), .CK(clk), .RN(rst_n), .Q(D1[95]) );
  DFFRHQX1 D1_reg_96_ ( .D(N5354), .CK(clk), .RN(rst_n), .Q(D1[96]) );
  DFFRHQX1 D1_reg_97_ ( .D(N5355), .CK(clk), .RN(rst_n), .Q(D1[97]) );
  DFFRHQX1 D1_reg_98_ ( .D(N5356), .CK(clk), .RN(rst_n), .Q(D1[98]) );
  DFFRHQX1 D1_reg_99_ ( .D(N5357), .CK(clk), .RN(rst_n), .Q(D1[99]) );
  DFFRHQX1 D1_reg_100_ ( .D(N5358), .CK(clk), .RN(rst_n), .Q(D1[100]) );
  DFFRHQX1 D1_reg_101_ ( .D(N5359), .CK(clk), .RN(rst_n), .Q(D1[101]) );
  DFFRHQX1 D1_reg_102_ ( .D(N5360), .CK(clk), .RN(rst_n), .Q(D1[102]) );
  DFFRHQX1 D1_reg_103_ ( .D(N5361), .CK(clk), .RN(rst_n), .Q(D1[103]) );
  DFFRHQX1 D1_reg_104_ ( .D(N5362), .CK(clk), .RN(rst_n), .Q(D1[104]) );
  DFFRHQX1 D1_reg_105_ ( .D(N5363), .CK(clk), .RN(rst_n), .Q(D1[105]) );
  DFFRHQX1 D1_reg_106_ ( .D(N5364), .CK(clk), .RN(rst_n), .Q(D1[106]) );
  DFFRHQX1 D1_reg_107_ ( .D(N5365), .CK(clk), .RN(rst_n), .Q(D1[107]) );
  DFFRHQX1 D1_reg_108_ ( .D(N5366), .CK(clk), .RN(rst_n), .Q(D1[108]) );
  DFFRHQX1 D1_reg_109_ ( .D(N5367), .CK(clk), .RN(rst_n), .Q(D1[109]) );
  DFFRHQX1 D1_reg_110_ ( .D(N5368), .CK(clk), .RN(rst_n), .Q(D1[110]) );
  DFFRHQX1 D1_reg_111_ ( .D(N5369), .CK(clk), .RN(rst_n), .Q(D1[111]) );
  DFFRHQX1 D1_reg_112_ ( .D(N5370), .CK(clk), .RN(rst_n), .Q(D1[112]) );
  DFFRHQX1 D1_reg_113_ ( .D(N5371), .CK(clk), .RN(rst_n), .Q(D1[113]) );
  DFFRHQX1 D1_reg_114_ ( .D(N5372), .CK(clk), .RN(rst_n), .Q(D1[114]) );
  DFFRHQX1 D1_reg_115_ ( .D(N5373), .CK(clk), .RN(rst_n), .Q(D1[115]) );
  DFFRHQX1 D1_reg_116_ ( .D(N5374), .CK(clk), .RN(rst_n), .Q(D1[116]) );
  DFFRHQX1 D1_reg_117_ ( .D(N5375), .CK(clk), .RN(rst_n), .Q(D1[117]) );
  DFFRHQX1 D1_reg_118_ ( .D(N5376), .CK(clk), .RN(rst_n), .Q(D1[118]) );
  DFFRHQX1 D1_reg_119_ ( .D(N5377), .CK(clk), .RN(rst_n), .Q(D1[119]) );
  DFFRHQX1 D1_reg_120_ ( .D(N5378), .CK(clk), .RN(rst_n), .Q(D1[120]) );
  DFFRHQX1 D1_reg_121_ ( .D(N5379), .CK(clk), .RN(rst_n), .Q(D1[121]) );
  DFFRHQX1 D1_reg_122_ ( .D(N5380), .CK(clk), .RN(rst_n), .Q(D1[122]) );
  DFFRHQX1 D1_reg_123_ ( .D(N5381), .CK(clk), .RN(rst_n), .Q(D1[123]) );
  DFFRHQX1 D1_reg_124_ ( .D(N5382), .CK(clk), .RN(rst_n), .Q(D1[124]) );
  DFFRHQX1 D1_reg_125_ ( .D(N5383), .CK(clk), .RN(rst_n), .Q(D1[125]) );
  DFFRHQX1 D1_reg_126_ ( .D(N5384), .CK(clk), .RN(rst_n), .Q(D1[126]) );
  DFFRHQX1 D3_reg_0_ ( .D(N5387), .CK(clk), .RN(rst_n), .Q(D3[0]) );
  DFFRHQX1 D3_reg_1_ ( .D(N5388), .CK(clk), .RN(rst_n), .Q(D3[1]) );
  DFFRHQX1 D3_reg_2_ ( .D(N5389), .CK(clk), .RN(rst_n), .Q(D3[2]) );
  DFFRHQX1 D3_reg_3_ ( .D(N5390), .CK(clk), .RN(rst_n), .Q(D3[3]) );
  DFFRHQX1 D3_reg_4_ ( .D(N5391), .CK(clk), .RN(rst_n), .Q(D3[4]) );
  DFFRHQX1 D3_reg_5_ ( .D(N5392), .CK(clk), .RN(rst_n), .Q(D3[5]) );
  DFFRHQX1 D3_reg_6_ ( .D(N5393), .CK(clk), .RN(rst_n), .Q(D3[6]) );
  DFFRHQX1 D3_reg_7_ ( .D(N5394), .CK(clk), .RN(rst_n), .Q(D3[7]) );
  DFFRHQX1 D3_reg_8_ ( .D(N5395), .CK(clk), .RN(rst_n), .Q(D3[8]) );
  DFFRHQX1 D3_reg_9_ ( .D(N5396), .CK(clk), .RN(rst_n), .Q(D3[9]) );
  DFFRHQX1 D3_reg_10_ ( .D(N5397), .CK(clk), .RN(rst_n), .Q(D3[10]) );
  DFFRHQX1 D3_reg_11_ ( .D(N5398), .CK(clk), .RN(rst_n), .Q(D3[11]) );
  DFFRHQX1 D3_reg_12_ ( .D(N5399), .CK(clk), .RN(rst_n), .Q(D3[12]) );
  DFFRHQX1 D3_reg_13_ ( .D(N5400), .CK(clk), .RN(rst_n), .Q(D3[13]) );
  DFFRHQX1 D3_reg_14_ ( .D(N5401), .CK(clk), .RN(rst_n), .Q(D3[14]) );
  DFFRHQX1 count78_reg_6_ ( .D(n3164), .CK(clk), .RN(rst_n), .Q(count78[6]) );
  DFFRHQX1 count68_reg_6_ ( .D(n3157), .CK(clk), .RN(rst_n), .Q(count68[6]) );
  DFFRHQX1 count28_reg_6_ ( .D(n3129), .CK(clk), .RN(rst_n), .Q(count28[6]) );
  DFFRHQX1 temp_i_mat_idx_reg_2_ ( .D(n2847), .CK(clk), .RN(rst_n), .Q(
        temp_i_mat_idx[2]) );
  DFFRHQX1 temp_i_mat_idx_reg_3_ ( .D(n2846), .CK(clk), .RN(rst_n), .Q(
        temp_i_mat_idx[3]) );
  DFFRHQX1 temp_i_mat_idx_reg_0_ ( .D(n2849), .CK(clk), .RN(rst_n), .Q(
        temp_i_mat_idx[0]) );
  DFFRHQX1 temp_i_mat_idx_reg_1_ ( .D(n2848), .CK(clk), .RN(rst_n), .Q(
        temp_i_mat_idx[1]) );
  DFFSHQX1 in_slut_reg ( .D(n4030), .CK(clk), .SN(rst_n), .Q(in_slut) );
  DFFRHQX1 count48_reg_6_ ( .D(n3143), .CK(clk), .RN(rst_n), .Q(count48[6]) );
  DFFRHQX1 count_state_idle_reg_5_ ( .D(n7198), .CK(clk), .RN(rst_n), .Q(
        count_state_idle[5]) );
  DFFRHQX1 A3_reg_6_ ( .D(N5151), .CK(clk), .RN(rst_n), .Q(A3[6]) );
  DFFRHQX1 count38_reg_6_ ( .D(n3136), .CK(clk), .RN(rst_n), .Q(count38[6]) );
  DFFRHQX1 count28_reg_5_ ( .D(n3130), .CK(clk), .RN(rst_n), .Q(count28[5]) );
  DFFRHQX1 count78_reg_5_ ( .D(n3165), .CK(clk), .RN(rst_n), .Q(count78[5]) );
  DFFRHQX1 count58_reg_6_ ( .D(n3150), .CK(clk), .RN(rst_n), .Q(count58[6]) );
  DFFRHQX1 count48_reg_5_ ( .D(n3144), .CK(clk), .RN(rst_n), .Q(count48[5]) );
  DFFRHQX1 count68_reg_5_ ( .D(n3158), .CK(clk), .RN(rst_n), .Q(count68[5]) );
  DFFRHQX1 count38_reg_5_ ( .D(n3137), .CK(clk), .RN(rst_n), .Q(count38[5]) );
  DFFRHQX1 count18_reg_6_ ( .D(n3122), .CK(clk), .RN(rst_n), .Q(count18[6]) );
  DFFRHQX1 reg_invalid2_signal_reg ( .D(n4001), .CK(clk), .RN(rst_n), .Q(
        reg_invalid2_signal) );
  DFFRHQX1 count58_reg_5_ ( .D(n3151), .CK(clk), .RN(rst_n), .Q(count58[5]) );
  DFFRHQX1 A3_reg_3_ ( .D(N5148), .CK(clk), .RN(rst_n), .Q(A3[3]) );
  DFFRHQX1 A3_reg_4_ ( .D(N5149), .CK(clk), .RN(rst_n), .Q(A3[4]) );
  DFFRHQX1 A3_reg_5_ ( .D(N5150), .CK(clk), .RN(rst_n), .Q(A3[5]) );
  DFFRHQX1 count08_reg_5_ ( .D(n3116), .CK(clk), .RN(rst_n), .Q(count08[5]) );
  DFFRHQX1 count38_reg_4_ ( .D(n3138), .CK(clk), .RN(rst_n), .Q(count38[4]) );
  DFFRHQX1 count48_reg_4_ ( .D(n3145), .CK(clk), .RN(rst_n), .Q(count48[4]) );
  DFFRHQX1 count58_reg_4_ ( .D(n3152), .CK(clk), .RN(rst_n), .Q(count58[4]) );
  DFFRHQX1 count68_reg_4_ ( .D(n3159), .CK(clk), .RN(rst_n), .Q(count68[4]) );
  DFFRHQX1 count28_reg_4_ ( .D(n3131), .CK(clk), .RN(rst_n), .Q(count28[4]) );
  DFFRHQX1 count78_reg_4_ ( .D(n3166), .CK(clk), .RN(rst_n), .Q(count78[4]) );
  DFFRHQX1 count_state_idle_reg_4_ ( .D(n7199), .CK(clk), .RN(rst_n), .Q(
        count_state_idle[4]) );
  DFFRHQX1 temp_w_mat_idx_reg_3_ ( .D(n2842), .CK(clk), .RN(rst_n), .Q(
        temp_w_mat_idx[3]) );
  DFFRHQX1 temp_w_mat_idx_reg_0_ ( .D(n2845), .CK(clk), .RN(rst_n), .Q(
        temp_w_mat_idx[0]) );
  DFFRHQX1 temp_w_mat_idx_reg_1_ ( .D(n2844), .CK(clk), .RN(rst_n), .Q(
        temp_w_mat_idx[1]) );
  DFFRHQX1 temp_w_mat_idx_reg_2_ ( .D(n2843), .CK(clk), .RN(rst_n), .Q(
        temp_w_mat_idx[2]) );
  DFFRHQX1 count08_reg_6_ ( .D(n3115), .CK(clk), .RN(rst_n), .Q(count08[6]) );
  DFFRHQX1 count08_reg_4_ ( .D(n3117), .CK(clk), .RN(rst_n), .Q(count08[4]) );
  DFFRHQX1 count18_reg_5_ ( .D(n3123), .CK(clk), .RN(rst_n), .Q(count18[5]) );
  DFFRHQX1 count18_reg_4_ ( .D(n3124), .CK(clk), .RN(rst_n), .Q(count18[4]) );
  DFFRHQX1 count_state_idle_reg_3_ ( .D(n7200), .CK(clk), .RN(rst_n), .Q(
        count_state_idle[3]) );
  DFFRHQX1 count38_reg_3_ ( .D(n3139), .CK(clk), .RN(rst_n), .Q(count38[3]) );
  DFFRHQX1 count48_reg_3_ ( .D(n3146), .CK(clk), .RN(rst_n), .Q(count48[3]) );
  DFFRHQX1 count58_reg_3_ ( .D(n3153), .CK(clk), .RN(rst_n), .Q(count58[3]) );
  DFFRHQX1 count_reg_15_ ( .D(n4011), .CK(clk), .RN(rst_n), .Q(count[15]) );
  DFFRHQX1 count18_reg_3_ ( .D(n3125), .CK(clk), .RN(rst_n), .Q(count18[3]) );
  DFFRHQX1 count68_reg_3_ ( .D(n3160), .CK(clk), .RN(rst_n), .Q(count68[3]) );
  DFFRHQX1 count08_reg_3_ ( .D(n3118), .CK(clk), .RN(rst_n), .Q(count08[3]) );
  DFFRHQX1 count28_reg_3_ ( .D(n3132), .CK(clk), .RN(rst_n), .Q(count28[3]) );
  DFFRHQX1 count78_reg_3_ ( .D(n3167), .CK(clk), .RN(rst_n), .Q(count78[3]) );
  DFFRHQX1 A3_reg_1_ ( .D(N5146), .CK(clk), .RN(rst_n), .Q(A3[1]) );
  DFFRHQX1 count1_reg_0_ ( .D(n7283), .CK(clk), .RN(rst_n), .Q(count1[0]) );
  DFFRHQX1 A3_reg_2_ ( .D(N5147), .CK(clk), .RN(rst_n), .Q(A3[2]) );
  DFFRHQX1 A3_reg_0_ ( .D(N5145), .CK(clk), .RN(rst_n), .Q(A3[0]) );
  DFFRHQX1 count_state_idle_reg_2_ ( .D(n7201), .CK(clk), .RN(rst_n), .Q(
        count_state_idle[2]) );
  DFFRHQX1 count1_reg_2_ ( .D(n3979), .CK(clk), .RN(rst_n), .Q(count1[2]) );
  DFFRHQX1 count_reg_14_ ( .D(n4012), .CK(clk), .RN(rst_n), .Q(count[14]) );
  DFFRHQX1 count58_reg_2_ ( .D(n3154), .CK(clk), .RN(rst_n), .Q(count58[2]) );
  DFFRHQX1 count08_reg_2_ ( .D(n3119), .CK(clk), .RN(rst_n), .Q(count08[2]) );
  DFFRHQX1 count28_reg_2_ ( .D(n3133), .CK(clk), .RN(rst_n), .Q(count28[2]) );
  DFFRHQX1 count48_reg_2_ ( .D(n3147), .CK(clk), .RN(rst_n), .Q(count48[2]) );
  DFFRHQX1 count78_reg_2_ ( .D(n3168), .CK(clk), .RN(rst_n), .Q(count78[2]) );
  DFFRHQX1 count38_reg_2_ ( .D(n3140), .CK(clk), .RN(rst_n), .Q(count38[2]) );
  DFFRHQX1 count18_reg_2_ ( .D(n3126), .CK(clk), .RN(rst_n), .Q(count18[2]) );
  DFFRHQX1 count68_reg_2_ ( .D(n3161), .CK(clk), .RN(rst_n), .Q(count68[2]) );
  DFFRHQX1 count1_reg_1_ ( .D(n3981), .CK(clk), .RN(rst_n), .Q(count1[1]) );
  DFFRHQX1 count08_reg_0_ ( .D(n3121), .CK(clk), .RN(rst_n), .Q(count08[0]) );
  DFFRHQX1 count18_reg_0_ ( .D(n3128), .CK(clk), .RN(rst_n), .Q(count18[0]) );
  DFFRHQX1 count_reg_12_ ( .D(n4014), .CK(clk), .RN(rst_n), .Q(count[12]) );
  DFFRHQX1 count58_reg_0_ ( .D(n3156), .CK(clk), .RN(rst_n), .Q(count58[0]) );
  DFFRHQX1 count28_reg_0_ ( .D(n3135), .CK(clk), .RN(rst_n), .Q(count28[0]) );
  DFFRHQX1 count78_reg_0_ ( .D(n3170), .CK(clk), .RN(rst_n), .Q(count78[0]) );
  DFFRHQX1 count48_reg_0_ ( .D(n3149), .CK(clk), .RN(rst_n), .Q(count48[0]) );
  DFFRHQX1 count38_reg_0_ ( .D(n3142), .CK(clk), .RN(rst_n), .Q(count38[0]) );
  DFFRHQX1 count68_reg_0_ ( .D(n3163), .CK(clk), .RN(rst_n), .Q(count68[0]) );
  DFFRHQXL reg_length00_reg_4_ ( .D(n3172), .CK(clk), .RN(rst_n), .Q(
        reg_length00[4]) );
  DFFRHQX1 count_state_idle_reg_1_ ( .D(n7202), .CK(clk), .RN(rst_n), .Q(
        count_state_idle[1]) );
  DFFRHQX1 count38_reg_1_ ( .D(n3141), .CK(clk), .RN(rst_n), .Q(count38[1]) );
  DFFRHQX1 count58_reg_1_ ( .D(n3155), .CK(clk), .RN(rst_n), .Q(count58[1]) );
  DFFRHQX1 count18_reg_1_ ( .D(n3127), .CK(clk), .RN(rst_n), .Q(count18[1]) );
  DFFRHQX1 count68_reg_1_ ( .D(n3162), .CK(clk), .RN(rst_n), .Q(count68[1]) );
  DFFRHQX1 count08_reg_1_ ( .D(n3120), .CK(clk), .RN(rst_n), .Q(count08[1]) );
  DFFRHQX1 count28_reg_1_ ( .D(n3134), .CK(clk), .RN(rst_n), .Q(count28[1]) );
  DFFRHQX1 count48_reg_1_ ( .D(n3148), .CK(clk), .RN(rst_n), .Q(count48[1]) );
  DFFRHQX1 count78_reg_1_ ( .D(n3169), .CK(clk), .RN(rst_n), .Q(count78[1]) );
  DFFRHQXL reg_length00_reg_5_ ( .D(n3171), .CK(clk), .RN(rst_n), .Q(
        reg_length00[5]) );
  DFFRHQXL reg_length00_reg_3_ ( .D(n3173), .CK(clk), .RN(rst_n), .Q(
        reg_length00[3]) );
  DFFRHQX1 count_reg_13_ ( .D(n4013), .CK(clk), .RN(rst_n), .Q(count[13]) );
  DFFRX1 count_state_idle_reg_0_ ( .D(n4002), .CK(clk), .RN(rst_n), .Q(
        count_state_idle[0]), .QN(n2858) );
  DFFRHQX1 count7_reg_2_ ( .D(n3568), .CK(clk), .RN(rst_n), .Q(count7[2]) );
  DFFRHQX1 count12_reg_0_ ( .D(n3294), .CK(clk), .RN(rst_n), .Q(count12[0]) );
  DFFRHQX1 count14_reg_0_ ( .D(n7268), .CK(clk), .RN(rst_n), .Q(count14[0]) );
  DFFRHQX1 count11_reg_2_ ( .D(n3348), .CK(clk), .RN(rst_n), .Q(count11[2]) );
  DFFRHQX1 count9_reg_2_ ( .D(n3458), .CK(clk), .RN(rst_n), .Q(count9[2]) );
  DFFRHQX1 count5_reg_2_ ( .D(n3678), .CK(clk), .RN(rst_n), .Q(count5[2]) );
  DFFRHQX1 count3_reg_2_ ( .D(n3788), .CK(clk), .RN(rst_n), .Q(count3[2]) );
  DFFRHQX1 count7_reg_0_ ( .D(n3569), .CK(clk), .RN(rst_n), .Q(count7[0]) );
  DFFRHQX1 count_reg_11_ ( .D(n4015), .CK(clk), .RN(rst_n), .Q(N5119) );
  DFFRHQX1 count8_reg_2_ ( .D(n3513), .CK(clk), .RN(rst_n), .Q(count8[2]) );
  DFFRHQX1 count2_reg_2_ ( .D(n3843), .CK(clk), .RN(rst_n), .Q(count2[2]) );
  DFFRHQX1 count5_reg_0_ ( .D(n3679), .CK(clk), .RN(rst_n), .Q(count5[0]) );
  DFFRHQX1 count6_reg_2_ ( .D(n3623), .CK(clk), .RN(rst_n), .Q(count6[2]) );
  DFFRHQX1 count10_reg_2_ ( .D(n3403), .CK(clk), .RN(rst_n), .Q(count10[2]) );
  DFFRHQX1 count11_reg_0_ ( .D(n3349), .CK(clk), .RN(rst_n), .Q(count11[0]) );
  DFFRHQX1 count9_reg_0_ ( .D(n3459), .CK(clk), .RN(rst_n), .Q(count9[0]) );
  DFFRHQX1 count11_reg_1_ ( .D(n3350), .CK(clk), .RN(rst_n), .Q(count11[1]) );
  DFFRHQX1 count3_reg_0_ ( .D(n3789), .CK(clk), .RN(rst_n), .Q(count3[0]) );
  DFFRHQX1 count4_reg_2_ ( .D(n3733), .CK(clk), .RN(rst_n), .Q(count4[2]) );
  DFFRHQX1 count12_reg_2_ ( .D(n3293), .CK(clk), .RN(rst_n), .Q(count12[2]) );
  DFFRHQX1 count9_reg_1_ ( .D(n3460), .CK(clk), .RN(rst_n), .Q(count9[1]) );
  DFFRHQX1 count7_reg_1_ ( .D(n3570), .CK(clk), .RN(rst_n), .Q(count7[1]) );
  DFFRHQX1 count2_reg_0_ ( .D(n3844), .CK(clk), .RN(rst_n), .Q(count2[0]) );
  DFFRHQX1 count14_reg_2_ ( .D(n3183), .CK(clk), .RN(rst_n), .Q(count14[2]) );
  DFFRHQX1 count5_reg_1_ ( .D(n3680), .CK(clk), .RN(rst_n), .Q(count5[1]) );
  DFFRHQX1 count8_reg_0_ ( .D(n3514), .CK(clk), .RN(rst_n), .Q(count8[0]) );
  DFFRHQX1 count3_reg_1_ ( .D(n3790), .CK(clk), .RN(rst_n), .Q(count3[1]) );
  DFFRHQX1 count6_reg_0_ ( .D(n3624), .CK(clk), .RN(rst_n), .Q(count6[0]) );
  DFFRX1 reg_length00_reg_0_ ( .D(n3176), .CK(clk), .RN(rst_n), .Q(n2839), 
        .QN(n4954) );
  DFFRHQX1 count10_reg_0_ ( .D(n3404), .CK(clk), .RN(rst_n), .Q(count10[0]) );
  DFFRHQX1 count4_reg_0_ ( .D(n3734), .CK(clk), .RN(rst_n), .Q(count4[0]) );
  DFFRHQX1 count13_reg_0_ ( .D(n3239), .CK(clk), .RN(rst_n), .Q(count13[0]) );
  DFFRHQX1 count10_reg_1_ ( .D(n3405), .CK(clk), .RN(rst_n), .Q(count10[1]) );
  DFFRHQX1 count8_reg_1_ ( .D(n3515), .CK(clk), .RN(rst_n), .Q(count8[1]) );
  DFFRHQX1 count14_reg_1_ ( .D(n3185), .CK(clk), .RN(rst_n), .Q(count14[1]) );
  DFFRHQX1 count2_reg_1_ ( .D(n3845), .CK(clk), .RN(rst_n), .Q(count2[1]) );
  DFFRHQX1 count13_reg_2_ ( .D(n3238), .CK(clk), .RN(rst_n), .Q(count13[2]) );
  DFFRHQX1 count6_reg_1_ ( .D(n3625), .CK(clk), .RN(rst_n), .Q(count6[1]) );
  DFFRHQX1 count4_reg_1_ ( .D(n3735), .CK(clk), .RN(rst_n), .Q(count4[1]) );
  DFFRHQX1 count12_reg_1_ ( .D(n3295), .CK(clk), .RN(rst_n), .Q(count12[1]) );
  DFFRHQX1 count13_reg_1_ ( .D(n3240), .CK(clk), .RN(rst_n), .Q(count13[1]) );
  DFFRHQX1 reg_length06_reg_5_ ( .D(n3626), .CK(clk), .RN(rst_n), .Q(
        reg_length06[5]) );
  DFFRHQX1 reg_length06_reg_3_ ( .D(n3628), .CK(clk), .RN(rst_n), .Q(
        reg_length06[3]) );
  DFFRHQX1 reg_length06_reg_4_ ( .D(n3627), .CK(clk), .RN(rst_n), .Q(
        reg_length06[4]) );
  DFFRHQX1 reg_length03_reg_1_ ( .D(n3795), .CK(clk), .RN(rst_n), .Q(
        reg_length03[1]) );
  DFFRHQXL y_out_sum12_reg_33_ ( .D(n3307), .CK(clk), .RN(rst_n), .Q(
        y_out_sum12[33]) );
  DFFRHQXL y_out_sum12_reg_32_ ( .D(n3308), .CK(clk), .RN(rst_n), .Q(
        y_out_sum12[32]) );
  DFFRHQX1 reg_length02_reg_1_ ( .D(n3850), .CK(clk), .RN(rst_n), .Q(
        reg_length02[1]) );
  DFFRHQX1 reg_length03_reg_2_ ( .D(n3794), .CK(clk), .RN(rst_n), .Q(
        reg_length03[2]) );
  DFFRHQX1 reg_length05_reg_1_ ( .D(n3685), .CK(clk), .RN(rst_n), .Q(
        reg_length05[1]) );
  DFFRHQXL y_out_sum9_reg_33_ ( .D(n3472), .CK(clk), .RN(rst_n), .Q(
        y_out_sum9[33]) );
  DFFRHQX1 reg_length02_reg_2_ ( .D(n3849), .CK(clk), .RN(rst_n), .Q(
        reg_length02[2]) );
  DFFRHQX1 reg_length014_reg_0_ ( .D(n3191), .CK(clk), .RN(rst_n), .Q(
        reg_length014[0]) );
  DFFRHQXL y_out_sum9_reg_32_ ( .D(n3473), .CK(clk), .RN(rst_n), .Q(
        y_out_sum9[32]) );
  DFFRHQXL y_out_sum13_reg_33_ ( .D(n3252), .CK(clk), .RN(rst_n), .Q(
        y_out_sum13[33]) );
  DFFRHQX1 reg_length01_reg_1_ ( .D(n3982), .CK(clk), .RN(rst_n), .Q(
        reg_length01[1]) );
  DFFRHQXL y_out_sum12_reg_37_ ( .D(n3303), .CK(clk), .RN(rst_n), .Q(
        y_out_sum12[37]) );
  DFFRHQX1 reg_length05_reg_2_ ( .D(n3684), .CK(clk), .RN(rst_n), .Q(
        reg_length05[2]) );
  DFFRHQXL y_out_sum12_reg_36_ ( .D(n3304), .CK(clk), .RN(rst_n), .Q(
        y_out_sum12[36]) );
  DFFRHQX1 reg_length011_reg_0_ ( .D(n3356), .CK(clk), .RN(rst_n), .Q(
        reg_length011[0]) );
  DFFRHQXL y_out_sum13_reg_32_ ( .D(n3253), .CK(clk), .RN(rst_n), .Q(
        y_out_sum13[32]) );
  DFFRHQX1 reg_length06_reg_0_ ( .D(n3631), .CK(clk), .RN(rst_n), .Q(
        reg_length06[0]) );
  DFFRHQX1 reg_length01_reg_2_ ( .D(n3983), .CK(clk), .RN(rst_n), .Q(
        reg_length01[2]) );
  DFFRHQXL y_out_sum9_reg_37_ ( .D(n3468), .CK(clk), .RN(rst_n), .Q(
        y_out_sum9[37]) );
  DFFRHQXL y_out_sum7_reg_33_ ( .D(n3582), .CK(clk), .RN(rst_n), .Q(
        y_out_sum7[33]) );
  DFFRHQX1 reg_length013_reg_3_ ( .D(n3243), .CK(clk), .RN(rst_n), .Q(
        reg_length013[3]) );
  DFFRHQXL y_out_sum7_reg_32_ ( .D(n3583), .CK(clk), .RN(rst_n), .Q(
        y_out_sum7[32]) );
  DFFRHQXL y_out_sum9_reg_36_ ( .D(n3469), .CK(clk), .RN(rst_n), .Q(
        y_out_sum9[36]) );
  DFFRHQX1 reg_length09_reg_0_ ( .D(n3466), .CK(clk), .RN(rst_n), .Q(
        reg_length09[0]) );
  DFFRHQXL y_out_sum13_reg_37_ ( .D(n3248), .CK(clk), .RN(rst_n), .Q(
        y_out_sum13[37]) );
  DFFRHQXL y_out_sum13_reg_36_ ( .D(n3249), .CK(clk), .RN(rst_n), .Q(
        y_out_sum13[36]) );
  DFFRHQX1 reg_length010_reg_0_ ( .D(n3411), .CK(clk), .RN(rst_n), .Q(
        reg_length010[0]) );
  DFFRHQX1 reg_length03_reg_3_ ( .D(n3793), .CK(clk), .RN(rst_n), .Q(
        reg_length03[3]) );
  DFFRHQX1 reg_length012_reg_0_ ( .D(n3301), .CK(clk), .RN(rst_n), .Q(
        reg_length012[0]) );
  DFFRHQX1 reg_length014_reg_3_ ( .D(n3188), .CK(clk), .RN(rst_n), .Q(
        reg_length014[3]) );
  DFFRHQXL y_out_sum7_reg_37_ ( .D(n3578), .CK(clk), .RN(rst_n), .Q(
        y_out_sum7[37]) );
  DFFRHQX1 reg_length07_reg_3_ ( .D(n3573), .CK(clk), .RN(rst_n), .Q(
        reg_length07[3]) );
  DFFRHQX1 reg_length013_reg_5_ ( .D(n3241), .CK(clk), .RN(rst_n), .Q(
        reg_length013[5]) );
  DFFRHQX1 reg_length011_reg_3_ ( .D(n3353), .CK(clk), .RN(rst_n), .Q(
        reg_length011[3]) );
  DFFRHQXL y_out_sum7_reg_36_ ( .D(n3579), .CK(clk), .RN(rst_n), .Q(
        y_out_sum7[36]) );
  DFFRHQX1 reg_length01_reg_3_ ( .D(n3984), .CK(clk), .RN(rst_n), .Q(
        reg_length01[3]) );
  DFFRHQX1 reg_length013_reg_4_ ( .D(n3242), .CK(clk), .RN(rst_n), .Q(
        reg_length013[4]) );
  DFFRHQX1 reg_length03_reg_5_ ( .D(n3791), .CK(clk), .RN(rst_n), .Q(
        reg_length03[5]) );
  DFFRHQX1 reg_length08_reg_0_ ( .D(n3521), .CK(clk), .RN(rst_n), .Q(
        reg_length08[0]) );
  DFFRHQX1 reg_length02_reg_3_ ( .D(n3848), .CK(clk), .RN(rst_n), .Q(
        reg_length02[3]) );
  DFFRHQX1 reg_length014_reg_5_ ( .D(n3186), .CK(clk), .RN(rst_n), .Q(
        reg_length014[5]) );
  DFFRHQX1 reg_length04_reg_1_ ( .D(n3740), .CK(clk), .RN(rst_n), .Q(
        reg_length04[1]) );
  DFFRHQX1 reg_length07_reg_5_ ( .D(n3571), .CK(clk), .RN(rst_n), .Q(
        reg_length07[5]) );
  DFFRHQX1 reg_length09_reg_3_ ( .D(n3463), .CK(clk), .RN(rst_n), .Q(
        reg_length09[3]) );
  DFFRHQX1 reg_length011_reg_5_ ( .D(n3351), .CK(clk), .RN(rst_n), .Q(
        reg_length011[5]) );
  DFFRHQX1 reg_length05_reg_3_ ( .D(n3683), .CK(clk), .RN(rst_n), .Q(
        reg_length05[3]) );
  DFFRHQX1 reg_length03_reg_4_ ( .D(n3792), .CK(clk), .RN(rst_n), .Q(
        reg_length03[4]) );
  DFFRHQX1 reg_length012_reg_3_ ( .D(n3298), .CK(clk), .RN(rst_n), .Q(
        reg_length012[3]) );
  DFFRHQX1 count_reg_10_ ( .D(n4016), .CK(clk), .RN(rst_n), .Q(N5118) );
  DFFRHQX1 reg_length014_reg_4_ ( .D(n3187), .CK(clk), .RN(rst_n), .Q(
        reg_length014[4]) );
  DFFRX1 reg_length014_reg_2_ ( .D(n3189), .CK(clk), .RN(rst_n), .QN(n4953) );
  DFFRHQX1 reg_length010_reg_3_ ( .D(n3408), .CK(clk), .RN(rst_n), .Q(
        reg_length010[3]) );
  DFFRHQX1 reg_length04_reg_2_ ( .D(n3739), .CK(clk), .RN(rst_n), .Q(
        reg_length04[2]) );
  DFFRHQX1 reg_length011_reg_4_ ( .D(n3352), .CK(clk), .RN(rst_n), .Q(
        reg_length011[4]) );
  DFFRHQX1 reg_length07_reg_4_ ( .D(n3572), .CK(clk), .RN(rst_n), .Q(
        reg_length07[4]) );
  DFFRHQX1 reg_length01_reg_5_ ( .D(n4010), .CK(clk), .RN(rst_n), .Q(
        reg_length01[5]) );
  DFFRX1 reg_length06_reg_2_ ( .D(n3629), .CK(clk), .RN(rst_n), .QN(n4948) );
  DFFRHQX1 reg_length02_reg_5_ ( .D(n3846), .CK(clk), .RN(rst_n), .Q(
        reg_length02[5]) );
  DFFRX1 reg_length014_reg_1_ ( .D(n3190), .CK(clk), .RN(rst_n), .QN(n4900) );
  DFFRHQX1 reg_length09_reg_5_ ( .D(n3461), .CK(clk), .RN(rst_n), .Q(
        reg_length09[5]) );
  DFFRHQX1 reg_length05_reg_5_ ( .D(n3681), .CK(clk), .RN(rst_n), .Q(
        reg_length05[5]) );
  DFFRHQX1 reg_length01_reg_4_ ( .D(n3985), .CK(clk), .RN(rst_n), .Q(
        reg_length01[4]) );
  DFFRHQX1 reg_length013_reg_0_ ( .D(n3246), .CK(clk), .RN(rst_n), .Q(
        reg_length013[0]) );
  DFFRHQX1 reg_length012_reg_5_ ( .D(n3296), .CK(clk), .RN(rst_n), .Q(
        reg_length012[5]) );
  DFFRHQX1 reg_length08_reg_3_ ( .D(n3518), .CK(clk), .RN(rst_n), .Q(
        reg_length08[3]) );
  DFFRHQX1 reg_length02_reg_4_ ( .D(n3847), .CK(clk), .RN(rst_n), .Q(
        reg_length02[4]) );
  DFFRX1 reg_length06_reg_1_ ( .D(n3630), .CK(clk), .RN(rst_n), .Q(n2821), 
        .QN(n4896) );
  DFFRHQX1 reg_length010_reg_5_ ( .D(n3406), .CK(clk), .RN(rst_n), .Q(
        reg_length010[5]) );
  DFFRX1 reg_length011_reg_2_ ( .D(n3354), .CK(clk), .RN(rst_n), .QN(n4951) );
  DFFRHQX1 reg_length09_reg_4_ ( .D(n3462), .CK(clk), .RN(rst_n), .Q(
        reg_length09[4]) );
  DFFRHQX1 reg_length05_reg_4_ ( .D(n3682), .CK(clk), .RN(rst_n), .Q(
        reg_length05[4]) );
  DFFRX1 reg_length09_reg_2_ ( .D(n3464), .CK(clk), .RN(rst_n), .QN(n4950) );
  DFFRHQX1 reg_length012_reg_4_ ( .D(n3297), .CK(clk), .RN(rst_n), .Q(
        reg_length012[4]) );
  DFFRHQX1 reg_length010_reg_4_ ( .D(n3407), .CK(clk), .RN(rst_n), .Q(
        reg_length010[4]) );
  DFFRX1 reg_length010_reg_2_ ( .D(n3409), .CK(clk), .RN(rst_n), .QN(n4949) );
  DFFRX1 reg_length011_reg_1_ ( .D(n3355), .CK(clk), .RN(rst_n), .QN(n4899) );
  DFFRHQX1 reg_length07_reg_0_ ( .D(n3576), .CK(clk), .RN(rst_n), .Q(
        reg_length07[0]) );
  DFFRHQXL y_out_sum0_reg_38_ ( .D(n3938), .CK(clk), .RN(rst_n), .Q(
        y_out_sum0[38]) );
  DFFRX1 reg_length09_reg_1_ ( .D(n3465), .CK(clk), .RN(rst_n), .QN(n4898) );
  DFFRHQX1 reg_length04_reg_3_ ( .D(n3738), .CK(clk), .RN(rst_n), .Q(
        reg_length04[3]) );
  DFFRHQXL y_out_sum0_reg_35_ ( .D(n3941), .CK(clk), .RN(rst_n), .Q(
        y_out_sum0[35]) );
  DFFRHQXL y_out_sum0_reg_39_ ( .D(n3977), .CK(clk), .RN(rst_n), .Q(
        y_out_sum0[39]) );
  DFFRHQXL y_out_sum0_reg_34_ ( .D(n3942), .CK(clk), .RN(rst_n), .Q(
        y_out_sum0[34]) );
  DFFRHQX1 reg_length08_reg_5_ ( .D(n3516), .CK(clk), .RN(rst_n), .Q(
        reg_length08[5]) );
  DFFRXL y_out_sum12_reg_35_ ( .D(n3305), .CK(clk), .RN(rst_n), .Q(
        y_out_sum12[35]), .QN(n6449) );
  DFFRX1 reg_length010_reg_1_ ( .D(n3410), .CK(clk), .RN(rst_n), .QN(n4897) );
  DFFRHQXL y_out_sum8_reg_33_ ( .D(n3527), .CK(clk), .RN(rst_n), .Q(
        y_out_sum8[33]) );
  DFFRHQXL y_out_sum8_reg_32_ ( .D(n3528), .CK(clk), .RN(rst_n), .Q(
        y_out_sum8[32]) );
  DFFRX1 reg_length012_reg_2_ ( .D(n3299), .CK(clk), .RN(rst_n), .QN(n4947) );
  DFFRHQX1 reg_length08_reg_4_ ( .D(n3517), .CK(clk), .RN(rst_n), .Q(
        reg_length08[4]) );
  DFFRXL y_out_sum9_reg_35_ ( .D(n3470), .CK(clk), .RN(rst_n), .Q(
        y_out_sum9[35]), .QN(n6613) );
  DFFRX1 reg_length012_reg_1_ ( .D(n3300), .CK(clk), .RN(rst_n), .QN(n4895) );
  DFFRHQX1 reg_length04_reg_5_ ( .D(n3736), .CK(clk), .RN(rst_n), .Q(
        reg_length04[5]) );
  DFFRHQXL y_out_sum8_reg_37_ ( .D(n3523), .CK(clk), .RN(rst_n), .Q(
        y_out_sum8[37]) );
  DFFRXL y_out_sum13_reg_35_ ( .D(n3250), .CK(clk), .RN(rst_n), .Q(
        y_out_sum13[35]), .QN(n6395) );
  DFFRHQXL y_out_sum0_reg_36_ ( .D(n3940), .CK(clk), .RN(rst_n), .Q(
        y_out_sum0[36]) );
  DFFRX1 reg_length03_reg_0_ ( .D(n3796), .CK(clk), .RN(rst_n), .Q(n2818) );
  DFFRHQXL y_out_sum0_reg_33_ ( .D(n3943), .CK(clk), .RN(rst_n), .Q(
        y_out_sum0[33]) );
  DFFRHQXL y_out_sum0_reg_37_ ( .D(n3939), .CK(clk), .RN(rst_n), .Q(
        y_out_sum0[37]) );
  DFFRHQXL y_out_sum0_reg_32_ ( .D(n3944), .CK(clk), .RN(rst_n), .Q(
        y_out_sum0[32]) );
  DFFRHQXL y_out_sum8_reg_36_ ( .D(n3524), .CK(clk), .RN(rst_n), .Q(
        y_out_sum8[36]) );
  DFFRHQXL y_out_sum10_reg_33_ ( .D(n3417), .CK(clk), .RN(rst_n), .Q(
        y_out_sum10[33]) );
  DFFRHQXL y_out_sum10_reg_37_ ( .D(n3413), .CK(clk), .RN(rst_n), .Q(
        y_out_sum10[37]) );
  DFFRX1 reg_length08_reg_2_ ( .D(n3519), .CK(clk), .RN(rst_n), .QN(n4946) );
  DFFRHQX1 reg_length04_reg_4_ ( .D(n3737), .CK(clk), .RN(rst_n), .Q(
        reg_length04[4]) );
  DFFRXL y_out_sum12_reg_34_ ( .D(n3306), .CK(clk), .RN(rst_n), .Q(
        y_out_sum12[34]), .QN(n6807) );
  DFFRXL y_out_sum7_reg_35_ ( .D(n3580), .CK(clk), .RN(rst_n), .Q(
        y_out_sum7[35]), .QN(n6725) );
  DFFRHQXL y_out_sum10_reg_36_ ( .D(n3414), .CK(clk), .RN(rst_n), .Q(
        y_out_sum10[36]) );
  DFFRX1 reg_length02_reg_0_ ( .D(n3851), .CK(clk), .RN(rst_n), .Q(n2817) );
  DFFRHQXL y_out_sum10_reg_32_ ( .D(n3418), .CK(clk), .RN(rst_n), .Q(
        y_out_sum10[32]) );
  DFFRX1 reg_length013_reg_2_ ( .D(n3244), .CK(clk), .RN(rst_n), .QN(n4945) );
  DFFRX1 reg_length08_reg_1_ ( .D(n3520), .CK(clk), .RN(rst_n), .QN(n4894) );
  DFFRX1 reg_length05_reg_0_ ( .D(n3686), .CK(clk), .RN(rst_n), .Q(n2820) );
  DFFRXL y_out_sum9_reg_34_ ( .D(n3471), .CK(clk), .RN(rst_n), .Q(
        y_out_sum9[34]), .QN(n6855) );
  DFFRX1 reg_length01_reg_0_ ( .D(n3986), .CK(clk), .RN(rst_n), .Q(n2816) );
  DFFRX1 reg_length013_reg_1_ ( .D(n3245), .CK(clk), .RN(rst_n), .Q(n2835), 
        .QN(n4893) );
  DFFRXL y_out_sum13_reg_34_ ( .D(n3251), .CK(clk), .RN(rst_n), .Q(
        y_out_sum13[34]), .QN(n6831) );
  DFFRXL y_out_sum12_reg_39_ ( .D(n3341), .CK(clk), .RN(rst_n), .Q(
        y_out_sum12[39]), .QN(n6496) );
  DFFRX1 reg_length07_reg_2_ ( .D(n3574), .CK(clk), .RN(rst_n), .QN(n4944) );
  DFFRXL y_out_sum12_reg_38_ ( .D(n3302), .CK(clk), .RN(rst_n), .Q(
        y_out_sum12[38]), .QN(n6811) );
  DFFRXL y_out_sum10_reg_38_ ( .D(n3412), .CK(clk), .RN(rst_n), .Q(
        y_out_sum10[38]), .QN(n6553) );
  DFFRXL y_out_sum10_reg_34_ ( .D(n3416), .CK(clk), .RN(rst_n), .Q(
        y_out_sum10[34]), .QN(n6559) );
  DFFRXL y_out_sum7_reg_34_ ( .D(n3581), .CK(clk), .RN(rst_n), .Q(
        y_out_sum7[34]), .QN(n6879) );
  DFFRHQXL y_out_sum3_reg_38_ ( .D(n3797), .CK(clk), .RN(rst_n), .Q(
        y_out_sum3[38]) );
  DFFRX1 reg_length07_reg_1_ ( .D(n3575), .CK(clk), .RN(rst_n), .Q(n2823), 
        .QN(n4892) );
  DFFRHQXL y_out_sum3_reg_35_ ( .D(n3800), .CK(clk), .RN(rst_n), .Q(
        y_out_sum3[35]) );
  DFFRHQXL y_out_sum3_reg_34_ ( .D(n3801), .CK(clk), .RN(rst_n), .Q(
        y_out_sum3[34]) );
  DFFRXL y_out_sum13_reg_39_ ( .D(n3286), .CK(clk), .RN(rst_n), .Q(
        y_out_sum13[39]), .QN(n6442) );
  DFFRXL y_out_sum13_reg_38_ ( .D(n3247), .CK(clk), .RN(rst_n), .Q(
        y_out_sum13[38]), .QN(n6835) );
  DFFRXL y_out_sum7_reg_39_ ( .D(n3616), .CK(clk), .RN(rst_n), .Q(
        y_out_sum7[39]), .QN(n6772) );
  DFFRHQXL y_out_sum14_reg_37_ ( .D(n3193), .CK(clk), .RN(rst_n), .Q(
        y_out_sum14[37]) );
  DFFRHQXL y_out_sum14_reg_33_ ( .D(n3197), .CK(clk), .RN(rst_n), .Q(
        y_out_sum14[33]) );
  DFFRXL y_out_sum7_reg_38_ ( .D(n3577), .CK(clk), .RN(rst_n), .Q(
        y_out_sum7[38]), .QN(n6883) );
  DFFRHQXL y_out_sum11_reg_33_ ( .D(n3362), .CK(clk), .RN(rst_n), .Q(
        y_out_sum11[33]) );
  DFFRXL y_out_sum10_reg_35_ ( .D(n3415), .CK(clk), .RN(rst_n), .Q(
        y_out_sum10[35]), .QN(n6557) );
  DFFRHQXL y_out_sum14_reg_36_ ( .D(n3194), .CK(clk), .RN(rst_n), .Q(
        y_out_sum14[36]) );
  DFFRHQXL y_out_sum11_reg_32_ ( .D(n3363), .CK(clk), .RN(rst_n), .Q(
        y_out_sum11[32]) );
  DFFRX1 reg_length04_reg_0_ ( .D(n3741), .CK(clk), .RN(rst_n), .Q(n2819) );
  DFFRHQXL y_out_sum14_reg_32_ ( .D(n3198), .CK(clk), .RN(rst_n), .Q(
        y_out_sum14[32]) );
  DFFRHQXL y_out_sum3_reg_33_ ( .D(n3802), .CK(clk), .RN(rst_n), .Q(
        y_out_sum3[33]) );
  DFFRHQXL y_out_sum3_reg_36_ ( .D(n3799), .CK(clk), .RN(rst_n), .Q(
        y_out_sum3[36]) );
  DFFRHQX1 y_out_sum12_reg_17_ ( .D(n3323), .CK(clk), .RN(rst_n), .Q(
        y_out_sum12[17]) );
  DFFRXL y_out_sum9_reg_38_ ( .D(n3467), .CK(clk), .RN(rst_n), .Q(
        y_out_sum9[38]), .QN(n6859) );
  DFFRHQXL y_out_sum3_reg_32_ ( .D(n3803), .CK(clk), .RN(rst_n), .Q(
        y_out_sum3[32]) );
  DFFRHQXL y_out_sum3_reg_37_ ( .D(n3798), .CK(clk), .RN(rst_n), .Q(
        y_out_sum3[37]) );
  DFFRHQXL y_out_sum11_reg_37_ ( .D(n3358), .CK(clk), .RN(rst_n), .Q(
        y_out_sum11[37]) );
  DFFRHQXL y_out_sum11_reg_36_ ( .D(n3359), .CK(clk), .RN(rst_n), .Q(
        y_out_sum11[36]) );
  DFFRHQX1 y_out_sum9_reg_17_ ( .D(n3488), .CK(clk), .RN(rst_n), .Q(
        y_out_sum9[17]) );
  DFFRXL y_out_sum10_reg_39_ ( .D(n3451), .CK(clk), .RN(rst_n), .Q(
        y_out_sum10[39]), .QN(n6606) );
  DFFRHQXL y_out_sum0_reg_29_ ( .D(n3947), .CK(clk), .RN(rst_n), .Q(
        y_out_sum0[29]) );
  DFFRHQXL y_out_sum0_reg_27_ ( .D(n3949), .CK(clk), .RN(rst_n), .Q(
        y_out_sum0[27]) );
  DFFRHQXL y_out_sum12_reg_29_ ( .D(n3311), .CK(clk), .RN(rst_n), .Q(
        y_out_sum12[29]) );
  DFFRXL y_out_sum8_reg_35_ ( .D(n3525), .CK(clk), .RN(rst_n), .Q(
        y_out_sum8[35]), .QN(n6669) );
  DFFRHQX1 y_out_sum0_reg_15_ ( .D(n3961), .CK(clk), .RN(rst_n), .Q(
        y_out_sum0[15]) );
  DFFRHQX1 y_out_sum13_reg_17_ ( .D(n3268), .CK(clk), .RN(rst_n), .Q(
        y_out_sum13[17]) );
  DFFRHQX1 y_out_sum10_reg_17_ ( .D(n3433), .CK(clk), .RN(rst_n), .Q(
        y_out_sum10[17]) );
  DFFRHQXL y_out_sum9_reg_29_ ( .D(n3476), .CK(clk), .RN(rst_n), .Q(
        y_out_sum9[29]) );
  DFFRHQXL y_out_sum0_reg_31_ ( .D(n3945), .CK(clk), .RN(rst_n), .Q(
        y_out_sum0[31]) );
  DFFRHQX1 y_out_sum7_reg_17_ ( .D(n3598), .CK(clk), .RN(rst_n), .Q(
        y_out_sum7[17]) );
  DFFRHQXL y_out_sum1_reg_38_ ( .D(n3898), .CK(clk), .RN(rst_n), .Q(
        y_out_sum1[38]) );
  DFFRHQX1 y_out_sum0_reg_17_ ( .D(n3959), .CK(clk), .RN(rst_n), .Q(
        y_out_sum0[17]) );
  DFFRHQXL y_out_sum12_reg_28_ ( .D(n3312), .CK(clk), .RN(rst_n), .Q(
        y_out_sum12[28]) );
  DFFRHQXL y_out_sum13_reg_29_ ( .D(n3256), .CK(clk), .RN(rst_n), .Q(
        y_out_sum13[29]) );
  DFFRHQX1 y_out_sum9_reg_16_ ( .D(n3489), .CK(clk), .RN(rst_n), .Q(
        y_out_sum9[16]) );
  DFFRHQX1 y_out_sum12_reg_21_ ( .D(n3319), .CK(clk), .RN(rst_n), .Q(
        y_out_sum12[21]) );
  DFFRHQXL y_out_sum1_reg_35_ ( .D(n3901), .CK(clk), .RN(rst_n), .Q(
        y_out_sum1[35]) );
  DFFRHQXL y_out_sum1_reg_34_ ( .D(n3902), .CK(clk), .RN(rst_n), .Q(
        y_out_sum1[34]) );
  DFFRHQXL y_out_sum0_reg_28_ ( .D(n3948), .CK(clk), .RN(rst_n), .Q(
        y_out_sum0[28]) );
  DFFRHQX1 y_out_sum0_reg_21_ ( .D(n3955), .CK(clk), .RN(rst_n), .Q(
        y_out_sum0[21]) );
  DFFRHQX1 y_out_sum0_reg_26_ ( .D(n3950), .CK(clk), .RN(rst_n), .Q(
        y_out_sum0[26]) );
  DFFRHQX1 y_out_sum0_reg_19_ ( .D(n3957), .CK(clk), .RN(rst_n), .Q(
        y_out_sum0[19]) );
  DFFRHQXL y_out_sum2_reg_38_ ( .D(n3852), .CK(clk), .RN(rst_n), .Q(
        y_out_sum2[38]) );
  DFFRHQXL y_out_sum10_reg_29_ ( .D(n3421), .CK(clk), .RN(rst_n), .Q(
        y_out_sum10[29]) );
  DFFRHQX1 y_out_sum0_reg_14_ ( .D(n3962), .CK(clk), .RN(rst_n), .Q(
        y_out_sum0[14]) );
  DFFRXL y_out_sum8_reg_34_ ( .D(n3526), .CK(clk), .RN(rst_n), .Q(
        y_out_sum8[34]), .QN(n6903) );
  DFFRHQXL y_out_sum9_reg_28_ ( .D(n3477), .CK(clk), .RN(rst_n), .Q(
        y_out_sum9[28]) );
  DFFRHQXL y_out_sum0_reg_30_ ( .D(n3946), .CK(clk), .RN(rst_n), .Q(
        y_out_sum0[30]) );
  DFFRHQX1 y_out_sum13_reg_16_ ( .D(n3269), .CK(clk), .RN(rst_n), .Q(
        y_out_sum13[16]) );
  DFFRHQX1 y_out_sum9_reg_21_ ( .D(n3484), .CK(clk), .RN(rst_n), .Q(
        y_out_sum9[21]) );
  DFFRHQXL y_out_sum2_reg_35_ ( .D(n3855), .CK(clk), .RN(rst_n), .Q(
        y_out_sum2[35]) );
  DFFRHQXL y_out_sum7_reg_29_ ( .D(n3586), .CK(clk), .RN(rst_n), .Q(
        y_out_sum7[29]) );
  DFFRXL y_out_sum12_reg_30_ ( .D(n3310), .CK(clk), .RN(rst_n), .Q(
        y_out_sum12[30]), .QN(n6456) );
  DFFRHQXL y_out_sum2_reg_33_ ( .D(n3857), .CK(clk), .RN(rst_n), .Q(
        y_out_sum2[33]) );
  DFFRHQXL y_out_sum13_reg_28_ ( .D(n3257), .CK(clk), .RN(rst_n), .Q(
        y_out_sum13[28]) );
  DFFRHQX1 y_out_sum12_reg_20_ ( .D(n3320), .CK(clk), .RN(rst_n), .Q(
        y_out_sum12[20]) );
  DFFRHQX1 y_out_sum7_reg_16_ ( .D(n3599), .CK(clk), .RN(rst_n), .Q(
        y_out_sum7[16]) );
  DFFRHQX1 y_out_sum10_reg_16_ ( .D(n3434), .CK(clk), .RN(rst_n), .Q(
        y_out_sum10[16]) );
  DFFRHQX1 y_out_sum13_reg_21_ ( .D(n3264), .CK(clk), .RN(rst_n), .Q(
        y_out_sum13[21]) );
  DFFRHQXL y_out_sum1_reg_33_ ( .D(n3903), .CK(clk), .RN(rst_n), .Q(
        y_out_sum1[33]) );
  DFFRHQX1 y_out_sum0_reg_16_ ( .D(n3960), .CK(clk), .RN(rst_n), .Q(
        y_out_sum0[16]) );
  DFFRHQXL y_out_sum2_reg_36_ ( .D(n3854), .CK(clk), .RN(rst_n), .Q(
        y_out_sum2[36]) );
  DFFRHQX1 reg_length12_reg_5_ ( .D(n3287), .CK(clk), .RN(rst_n), .Q(
        reg_length12[5]) );
  DFFRHQXL y_out_sum7_reg_28_ ( .D(n3587), .CK(clk), .RN(rst_n), .Q(
        y_out_sum7[28]) );
  DFFRHQXL y_out_sum10_reg_28_ ( .D(n3422), .CK(clk), .RN(rst_n), .Q(
        y_out_sum10[28]) );
  DFFRHQXL y_out_sum1_reg_36_ ( .D(n3900), .CK(clk), .RN(rst_n), .Q(
        y_out_sum1[36]) );
  DFFRHQX1 y_out_sum9_reg_25_ ( .D(n3480), .CK(clk), .RN(rst_n), .Q(
        y_out_sum9[25]) );
  DFFRHQX1 y_out_sum10_reg_21_ ( .D(n3429), .CK(clk), .RN(rst_n), .Q(
        y_out_sum10[21]) );
  DFFRHQXL y_out_sum2_reg_34_ ( .D(n3856), .CK(clk), .RN(rst_n), .Q(
        y_out_sum2[34]) );
  DFFRHQX1 y_out_sum0_reg_20_ ( .D(n3956), .CK(clk), .RN(rst_n), .Q(
        y_out_sum0[20]) );
  DFFRHQXL y_out_sum1_reg_32_ ( .D(n3904), .CK(clk), .RN(rst_n), .Q(
        y_out_sum1[32]) );
  DFFRHQXL y_out_sum1_reg_37_ ( .D(n3899), .CK(clk), .RN(rst_n), .Q(
        y_out_sum1[37]) );
  DFFRHQX1 y_out_sum0_reg_18_ ( .D(n3958), .CK(clk), .RN(rst_n), .Q(
        y_out_sum0[18]) );
  DFFRHQX1 y_out_sum7_reg_21_ ( .D(n3594), .CK(clk), .RN(rst_n), .Q(
        y_out_sum7[21]) );
  DFFRHQX1 y_out_sum9_reg_20_ ( .D(n3485), .CK(clk), .RN(rst_n), .Q(
        y_out_sum9[20]) );
  DFFRXL y_out_sum8_reg_39_ ( .D(n3561), .CK(clk), .RN(rst_n), .Q(
        y_out_sum8[39]), .QN(n6717) );
  DFFRXL y_out_sum9_reg_30_ ( .D(n3475), .CK(clk), .RN(rst_n), .Q(
        y_out_sum9[30]), .QN(n6620) );
  DFFRXL y_out_sum8_reg_38_ ( .D(n3522), .CK(clk), .RN(rst_n), .Q(
        y_out_sum8[38]), .QN(n6907) );
  DFFRHQXL y_out_sum2_reg_32_ ( .D(n3858), .CK(clk), .RN(rst_n), .Q(
        y_out_sum2[32]) );
  DFFRHQX1 y_out_sum13_reg_25_ ( .D(n3260), .CK(clk), .RN(rst_n), .Q(
        y_out_sum13[25]) );
  DFFRHQX1 reg_length9_reg_5_ ( .D(n3452), .CK(clk), .RN(rst_n), .Q(
        reg_length9[5]) );
  DFFRX1 y_out_sum12_reg_22_ ( .D(n3318), .CK(clk), .RN(rst_n), .Q(
        y_out_sum12[22]), .QN(n4963) );
  DFFRHQX1 y_out_sum1_reg_39_ ( .D(n3937), .CK(clk), .RN(rst_n), .Q(
        y_out_sum1[39]) );
  DFFRXL y_out_sum13_reg_30_ ( .D(n3255), .CK(clk), .RN(rst_n), .Q(
        y_out_sum13[30]), .QN(n6402) );
  DFFRHQX1 y_out_sum9_reg_24_ ( .D(n3481), .CK(clk), .RN(rst_n), .Q(
        y_out_sum9[24]) );
  DFFRHQX1 y_out_sum13_reg_20_ ( .D(n3265), .CK(clk), .RN(rst_n), .Q(
        y_out_sum13[20]) );
  DFFRXL y_out_sum12_reg_31_ ( .D(n3309), .CK(clk), .RN(rst_n), .Q(
        y_out_sum12[31]), .QN(n6454) );
  DFFRXL y_out_sum10_reg_30_ ( .D(n3420), .CK(clk), .RN(rst_n), .Q(
        y_out_sum10[30]), .QN(n6565) );
  DFFRHQX1 y_out_sum13_reg_24_ ( .D(n3261), .CK(clk), .RN(rst_n), .Q(
        y_out_sum13[24]) );
  DFFRHQX1 y_out_sum10_reg_20_ ( .D(n3430), .CK(clk), .RN(rst_n), .Q(
        y_out_sum10[20]) );
  DFFRHQX1 y_out_sum12_reg_16_ ( .D(n3324), .CK(clk), .RN(rst_n), .Q(
        y_out_sum12[16]) );
  DFFRHQX1 y_out_sum7_reg_20_ ( .D(n3595), .CK(clk), .RN(rst_n), .Q(
        y_out_sum7[20]) );
  DFFRXL y_out_sum7_reg_30_ ( .D(n3585), .CK(clk), .RN(rst_n), .Q(
        y_out_sum7[30]), .QN(n6732) );
  DFFRHQXL y_out_sum3_reg_29_ ( .D(n3806), .CK(clk), .RN(rst_n), .Q(
        y_out_sum3[29]) );
  DFFRHQXL y_out_sum2_reg_37_ ( .D(n3853), .CK(clk), .RN(rst_n), .Q(
        y_out_sum2[37]) );
  DFFRHQX1 y_out_sum13_reg_13_ ( .D(n3272), .CK(clk), .RN(rst_n), .Q(
        y_out_sum13[13]) );
  DFFRX1 y_out_sum13_reg_22_ ( .D(n3263), .CK(clk), .RN(rst_n), .Q(
        y_out_sum13[22]), .QN(n4965) );
  DFFRHQX1 reg_length12_reg_4_ ( .D(n3288), .CK(clk), .RN(rst_n), .Q(
        reg_length12[4]) );
  DFFRHQXL y_out_sum3_reg_27_ ( .D(n3808), .CK(clk), .RN(rst_n), .Q(
        y_out_sum3[27]) );
  DFFRXL y_out_sum9_reg_31_ ( .D(n3474), .CK(clk), .RN(rst_n), .Q(
        y_out_sum9[31]), .QN(n6618) );
  DFFRHQX1 y_out_sum3_reg_15_ ( .D(n3820), .CK(clk), .RN(rst_n), .Q(
        y_out_sum3[15]) );
  DFFRHQX1 y_out_sum9_reg_13_ ( .D(n3492), .CK(clk), .RN(rst_n), .Q(
        y_out_sum9[13]) );
  DFFRHQXL y_out_sum3_reg_31_ ( .D(n3804), .CK(clk), .RN(rst_n), .Q(
        y_out_sum3[31]) );
  DFFRHQX1 y_out_sum3_reg_25_ ( .D(n3810), .CK(clk), .RN(rst_n), .Q(
        y_out_sum3[25]) );
  DFFRHQXL y_out_sum5_reg_38_ ( .D(n3687), .CK(clk), .RN(rst_n), .Q(
        y_out_sum5[38]) );
  DFFRHQX1 reg_length9_reg_4_ ( .D(n3453), .CK(clk), .RN(rst_n), .Q(
        reg_length9[4]) );
  DFFRXL y_out_sum13_reg_31_ ( .D(n3254), .CK(clk), .RN(rst_n), .Q(
        y_out_sum13[31]), .QN(n6400) );
  DFFRXL y_out_sum11_reg_35_ ( .D(n3360), .CK(clk), .RN(rst_n), .Q(
        y_out_sum11[35]), .QN(n6502) );
  DFFRHQX1 y_out_sum3_reg_13_ ( .D(n3822), .CK(clk), .RN(rst_n), .Q(
        y_out_sum3[13]) );
  DFFRXL y_out_sum12_reg_27_ ( .D(n3313), .CK(clk), .RN(rst_n), .Q(
        y_out_sum12[27]), .QN(n6460) );
  DFFRHQXL y_out_sum5_reg_35_ ( .D(n3690), .CK(clk), .RN(rst_n), .Q(
        y_out_sum5[35]) );
  DFFRX1 y_out_sum7_reg_22_ ( .D(n3593), .CK(clk), .RN(rst_n), .Q(
        y_out_sum7[22]), .QN(n4961) );
  DFFRHQXL y_out_sum5_reg_34_ ( .D(n3691), .CK(clk), .RN(rst_n), .Q(
        y_out_sum5[34]) );
  DFFRHQX1 y_out_sum0_reg_13_ ( .D(n3963), .CK(clk), .RN(rst_n), .Q(
        y_out_sum0[13]) );
  DFFRXL y_out_sum10_reg_31_ ( .D(n3419), .CK(clk), .RN(rst_n), .Q(
        y_out_sum10[31]), .QN(n6563) );
  DFFRX1 y_out_sum12_reg_23_ ( .D(n3317), .CK(clk), .RN(rst_n), .Q(
        y_out_sum12[23]), .QN(n4956) );
  DFFRHQX1 y_out_sum3_reg_14_ ( .D(n3821), .CK(clk), .RN(rst_n), .Q(
        y_out_sum3[14]) );
  DFFRHQX1 count_reg_9_ ( .D(n4017), .CK(clk), .RN(rst_n), .Q(N5062) );
  DFFRXL y_out_sum9_reg_27_ ( .D(n3478), .CK(clk), .RN(rst_n), .Q(
        y_out_sum9[27]), .QN(n6624) );
  DFFRXL y_out_sum14_reg_35_ ( .D(n3195), .CK(clk), .RN(rst_n), .Q(
        y_out_sum14[35]), .QN(n6341) );
  DFFRHQX1 y_out_sum10_reg_13_ ( .D(n3437), .CK(clk), .RN(rst_n), .Q(
        y_out_sum10[13]) );
  DFFRX1 y_out_sum10_reg_26_ ( .D(n3424), .CK(clk), .RN(rst_n), .Q(
        y_out_sum10[26]), .QN(n4958) );
  DFFRHQX1 reg_length13_reg_5_ ( .D(n3232), .CK(clk), .RN(rst_n), .Q(
        reg_length13[5]) );
  DFFRHQX1 y_out_sum8_reg_17_ ( .D(n3543), .CK(clk), .RN(rst_n), .Q(
        y_out_sum8[17]) );
  DFFRHQX1 count_reg_8_ ( .D(n4018), .CK(clk), .RN(rst_n), .Q(N5061) );
  DFFRXL y_out_sum7_reg_31_ ( .D(n3584), .CK(clk), .RN(rst_n), .Q(
        y_out_sum7[31]), .QN(n6730) );
  DFFRHQX1 reg_length3_reg_5_ ( .D(n3782), .CK(clk), .RN(rst_n), .Q(
        reg_length3[5]) );
  DFFRHQX1 y_out_sum3_reg_17_ ( .D(n3818), .CK(clk), .RN(rst_n), .Q(
        y_out_sum3[17]) );
  DFFRX1 y_out_sum7_reg_26_ ( .D(n3589), .CK(clk), .RN(rst_n), .Q(
        y_out_sum7[26]), .QN(n4959) );
  DFFRHQX1 y_out_sum7_reg_13_ ( .D(n3602), .CK(clk), .RN(rst_n), .Q(
        y_out_sum7[13]) );
  DFFRHQXL y_out_sum3_reg_30_ ( .D(n3805), .CK(clk), .RN(rst_n), .Q(
        y_out_sum3[30]) );
  DFFRXL y_out_sum13_reg_27_ ( .D(n3258), .CK(clk), .RN(rst_n), .Q(
        y_out_sum13[27]), .QN(n6406) );
  DFFRHQXL y_out_sum5_reg_33_ ( .D(n3692), .CK(clk), .RN(rst_n), .Q(
        y_out_sum5[33]) );
  DFFRHQX1 y_out_sum3_reg_21_ ( .D(n3814), .CK(clk), .RN(rst_n), .Q(
        y_out_sum3[21]) );
  DFFRXL y_out_sum14_reg_39_ ( .D(n3231), .CK(clk), .RN(rst_n), .Q(
        y_out_sum14[39]), .QN(n6388) );
  DFFRXL y_out_sum10_reg_27_ ( .D(n3423), .CK(clk), .RN(rst_n), .Q(
        y_out_sum10[27]), .QN(n6569) );
  DFFRXL y_out_sum14_reg_38_ ( .D(n3192), .CK(clk), .RN(rst_n), .Q(
        y_out_sum14[38]), .QN(n6951) );
  DFFRHQXL y_out_sum3_reg_28_ ( .D(n3807), .CK(clk), .RN(rst_n), .Q(
        y_out_sum3[28]) );
  DFFRX1 y_out_sum13_reg_23_ ( .D(n3262), .CK(clk), .RN(rst_n), .Q(
        y_out_sum13[23]), .QN(n4955) );
  DFFRHQXL y_out_sum5_reg_36_ ( .D(n3689), .CK(clk), .RN(rst_n), .Q(
        y_out_sum5[36]) );
  DFFRHQX1 y_out_sum3_reg_24_ ( .D(n3811), .CK(clk), .RN(rst_n), .Q(
        y_out_sum3[24]) );
  DFFRXL y_out_sum11_reg_34_ ( .D(n3361), .CK(clk), .RN(rst_n), .Q(
        y_out_sum11[34]), .QN(n6927) );
  DFFRHQXL y_out_sum8_reg_29_ ( .D(n3531), .CK(clk), .RN(rst_n), .Q(
        y_out_sum8[29]) );
  DFFRHQXL y_out_sum5_reg_32_ ( .D(n3693), .CK(clk), .RN(rst_n), .Q(
        y_out_sum5[32]) );
  DFFRHQXL y_out_sum5_reg_37_ ( .D(n3688), .CK(clk), .RN(rst_n), .Q(
        y_out_sum5[37]) );
  DFFRHQXL y_out_sum3_reg_26_ ( .D(n3809), .CK(clk), .RN(rst_n), .Q(
        y_out_sum3[26]) );
  DFFRXL y_out_sum7_reg_27_ ( .D(n3588), .CK(clk), .RN(rst_n), .Q(
        y_out_sum7[27]), .QN(n6736) );
  DFFRHQX1 reg_length13_reg_4_ ( .D(n3233), .CK(clk), .RN(rst_n), .Q(
        reg_length13[4]) );
  DFFRHQX1 y_out_sum3_reg_19_ ( .D(n3816), .CK(clk), .RN(rst_n), .Q(
        y_out_sum3[19]) );
  DFFRXL y_out_sum14_reg_34_ ( .D(n3196), .CK(clk), .RN(rst_n), .Q(
        y_out_sum14[34]), .QN(n6955) );
  DFFRHQX1 y_out_sum5_reg_39_ ( .D(n3726), .CK(clk), .RN(rst_n), .Q(
        y_out_sum5[39]) );
  DFFRX1 y_out_sum12_reg_18_ ( .D(n3322), .CK(clk), .RN(rst_n), .Q(
        y_out_sum12[18]), .QN(n4941) );
  DFFRHQX1 y_out_sum1_reg_13_ ( .D(n3923), .CK(clk), .RN(rst_n), .Q(
        y_out_sum1[13]) );
  DFFRHQX1 y_out_sum8_reg_16_ ( .D(n3544), .CK(clk), .RN(rst_n), .Q(
        y_out_sum8[16]) );
  DFFRHQX1 y_out_sum2_reg_39_ ( .D(n3891), .CK(clk), .RN(rst_n), .Q(
        y_out_sum2[39]) );
  DFFRHQX1 reg_length7_reg_4_ ( .D(n3563), .CK(clk), .RN(rst_n), .Q(
        reg_length7[4]) );
  DFFRHQX1 y_out_sum3_reg_16_ ( .D(n3819), .CK(clk), .RN(rst_n), .Q(
        y_out_sum3[16]) );
  DFFRHQX1 reg_length1_reg_5_ ( .D(n3892), .CK(clk), .RN(rst_n), .Q(
        reg_length1[5]) );
  DFFRHQX1 y_out_sum3_reg_18_ ( .D(n3817), .CK(clk), .RN(rst_n), .Q(
        y_out_sum3[18]) );
  DFFRHQX1 reg_length10_reg_4_ ( .D(n3398), .CK(clk), .RN(rst_n), .Q(
        reg_length10[4]) );
  DFFRHQXL y_out_sum8_reg_28_ ( .D(n3532), .CK(clk), .RN(rst_n), .Q(
        y_out_sum8[28]) );
  DFFRHQX1 y_out_sum8_reg_21_ ( .D(n3539), .CK(clk), .RN(rst_n), .Q(
        y_out_sum8[21]) );
  DFFRXL y_out_sum11_reg_39_ ( .D(n3396), .CK(clk), .RN(rst_n), .Q(
        y_out_sum11[39]), .QN(n6550) );
  DFFRHQX1 reg_length10_reg_5_ ( .D(n3397), .CK(clk), .RN(rst_n), .Q(
        reg_length10[5]) );
  DFFRXL y_out_sum11_reg_38_ ( .D(n3357), .CK(clk), .RN(rst_n), .Q(
        y_out_sum11[38]), .QN(n6931) );
  DFFRHQXL y_out_sum1_reg_29_ ( .D(n3907), .CK(clk), .RN(rst_n), .Q(
        y_out_sum1[29]) );
  DFFRX1 y_out_sum12_reg_19_ ( .D(n3321), .CK(clk), .RN(rst_n), .Q(
        y_out_sum12[19]), .QN(n4889) );
  DFFRX1 y_out_sum9_reg_18_ ( .D(n3487), .CK(clk), .RN(rst_n), .Q(
        y_out_sum9[18]), .QN(n4935) );
  DFFRX1 y_out_sum13_reg_18_ ( .D(n3267), .CK(clk), .RN(rst_n), .Q(
        y_out_sum13[18]), .QN(n4936) );
  DFFRHQX1 y_out_sum3_reg_20_ ( .D(n3815), .CK(clk), .RN(rst_n), .Q(
        y_out_sum3[20]) );
  DFFRHQXL y_out_sum6_reg_38_ ( .D(n3632), .CK(clk), .RN(rst_n), .Q(
        y_out_sum6[38]) );
  DFFRHQX1 y_out_sum1_reg_15_ ( .D(n3921), .CK(clk), .RN(rst_n), .Q(
        y_out_sum1[15]) );
  DFFRHQXL y_out_sum1_reg_31_ ( .D(n3905), .CK(clk), .RN(rst_n), .Q(
        y_out_sum1[31]) );
  DFFRHQX1 y_out_sum1_reg_25_ ( .D(n3911), .CK(clk), .RN(rst_n), .Q(
        y_out_sum1[25]) );
  DFFRHQX1 y_out_sum8_reg_25_ ( .D(n3535), .CK(clk), .RN(rst_n), .Q(
        y_out_sum8[25]) );
  DFFRX1 y_out_sum10_reg_18_ ( .D(n3432), .CK(clk), .RN(rst_n), .Q(
        y_out_sum10[18]), .QN(n4925) );
  DFFRHQXL y_out_sum1_reg_27_ ( .D(n3909), .CK(clk), .RN(rst_n), .Q(
        y_out_sum1[27]) );
  DFFRHQXL y_out_sum6_reg_35_ ( .D(n3635), .CK(clk), .RN(rst_n), .Q(
        y_out_sum6[35]) );
  DFFRXL y_out_sum8_reg_30_ ( .D(n3530), .CK(clk), .RN(rst_n), .Q(
        y_out_sum8[30]), .QN(n6676) );
  DFFRHQXL y_out_sum6_reg_34_ ( .D(n3636), .CK(clk), .RN(rst_n), .Q(
        y_out_sum6[34]) );
  DFFRHQX1 y_out_sum12_reg_13_ ( .D(n3327), .CK(clk), .RN(rst_n), .Q(
        y_out_sum12[13]) );
  DFFRX1 y_out_sum7_reg_18_ ( .D(n3597), .CK(clk), .RN(rst_n), .Q(
        y_out_sum7[18]), .QN(n4924) );
  DFFRHQX1 y_out_sum8_reg_20_ ( .D(n3540), .CK(clk), .RN(rst_n), .Q(
        y_out_sum8[20]) );
  DFFRX1 y_out_sum9_reg_19_ ( .D(n3486), .CK(clk), .RN(rst_n), .Q(
        y_out_sum9[19]), .QN(n4882) );
  DFFRHQX1 y_out_sum1_reg_14_ ( .D(n3922), .CK(clk), .RN(rst_n), .Q(
        y_out_sum1[14]) );
  DFFRHQX1 y_out_sum2_reg_13_ ( .D(n3877), .CK(clk), .RN(rst_n), .Q(
        y_out_sum2[13]) );
  DFFRX1 y_out_sum13_reg_19_ ( .D(n3266), .CK(clk), .RN(rst_n), .Q(
        y_out_sum13[19]), .QN(n4884) );
  DFFRHQX1 reg_length2_reg_5_ ( .D(n3837), .CK(clk), .RN(rst_n), .Q(
        reg_length2[5]) );
  DFFRHQX1 y_out_sum8_reg_24_ ( .D(n3536), .CK(clk), .RN(rst_n), .Q(
        y_out_sum8[24]) );
  DFFRHQX1 reg_length3_reg_4_ ( .D(n3783), .CK(clk), .RN(rst_n), .Q(
        reg_length3[4]) );
  DFFRHQX1 y_out_sum1_reg_17_ ( .D(n3919), .CK(clk), .RN(rst_n), .Q(
        y_out_sum1[17]) );
  DFFRHQXL y_out_sum4_reg_38_ ( .D(n3742), .CK(clk), .RN(rst_n), .Q(
        y_out_sum4[38]) );
  DFFRX1 y_out_sum10_reg_19_ ( .D(n3431), .CK(clk), .RN(rst_n), .Q(
        y_out_sum10[19]), .QN(n4873) );
  DFFRHQX1 y_out_sum8_reg_13_ ( .D(n3547), .CK(clk), .RN(rst_n), .Q(
        y_out_sum8[13]) );
  DFFRHQXL y_out_sum1_reg_30_ ( .D(n3906), .CK(clk), .RN(rst_n), .Q(
        y_out_sum1[30]) );
  DFFRHQXL y_out_sum4_reg_35_ ( .D(n3745), .CK(clk), .RN(rst_n), .Q(
        y_out_sum4[35]) );
  DFFRX1 y_out_sum7_reg_19_ ( .D(n3596), .CK(clk), .RN(rst_n), .Q(
        y_out_sum7[19]), .QN(n4872) );
  DFFRHQXL y_out_sum1_reg_28_ ( .D(n3908), .CK(clk), .RN(rst_n), .Q(
        y_out_sum1[28]) );
  DFFRHQX1 y_out_sum14_reg_17_ ( .D(n3213), .CK(clk), .RN(rst_n), .Q(
        y_out_sum14[17]) );
  DFFRX1 y_out_sum8_reg_22_ ( .D(n3538), .CK(clk), .RN(rst_n), .Q(
        y_out_sum8[22]), .QN(n4964) );
  DFFRHQXL y_out_sum4_reg_34_ ( .D(n3746), .CK(clk), .RN(rst_n), .Q(
        y_out_sum4[34]) );
  DFFRHQX1 y_out_sum1_reg_21_ ( .D(n3915), .CK(clk), .RN(rst_n), .Q(
        y_out_sum1[21]) );
  DFFRHQX1 y_out_sum2_reg_14_ ( .D(n3876), .CK(clk), .RN(rst_n), .Q(
        y_out_sum2[14]) );
  DFFRHQXL y_out_sum2_reg_29_ ( .D(n3861), .CK(clk), .RN(rst_n), .Q(
        y_out_sum2[29]) );
  DFFRHQXL y_out_sum6_reg_36_ ( .D(n3634), .CK(clk), .RN(rst_n), .Q(
        y_out_sum6[36]) );
  DFFRHQXL y_out_sum6_reg_33_ ( .D(n3637), .CK(clk), .RN(rst_n), .Q(
        y_out_sum6[33]) );
  DFFRHQXL y_out_sum2_reg_27_ ( .D(n3863), .CK(clk), .RN(rst_n), .Q(
        y_out_sum2[27]) );
  DFFRHQX1 y_out_sum1_reg_24_ ( .D(n3912), .CK(clk), .RN(rst_n), .Q(
        y_out_sum1[24]) );
  DFFRXL y_out_sum8_reg_31_ ( .D(n3529), .CK(clk), .RN(rst_n), .Q(
        y_out_sum8[31]), .QN(n6674) );
  DFFRHQXL y_out_sum6_reg_32_ ( .D(n3638), .CK(clk), .RN(rst_n), .Q(
        y_out_sum6[32]) );
  DFFRHQX1 y_out_sum0_reg_12_ ( .D(n3964), .CK(clk), .RN(rst_n), .Q(
        y_out_sum0[12]) );
  DFFRHQXL y_out_sum6_reg_37_ ( .D(n3633), .CK(clk), .RN(rst_n), .Q(
        y_out_sum6[37]) );
  DFFRHQX1 y_out_sum11_reg_17_ ( .D(n3378), .CK(clk), .RN(rst_n), .Q(
        y_out_sum11[17]) );
  DFFRHQX1 y_out_sum2_reg_17_ ( .D(n3873), .CK(clk), .RN(rst_n), .Q(
        y_out_sum2[17]) );
  DFFRX1 reg_length7_reg_5_ ( .D(n3562), .CK(clk), .RN(rst_n), .Q(
        reg_length7[5]), .QN(n5027) );
  DFFRHQX1 y_out_sum9_reg_12_ ( .D(n3493), .CK(clk), .RN(rst_n), .Q(
        y_out_sum9[12]) );
  DFFRHQX1 reg_length8_reg_5_ ( .D(n3507), .CK(clk), .RN(rst_n), .Q(
        reg_length8[5]) );
  DFFRHQXL y_out_sum2_reg_30_ ( .D(n3860), .CK(clk), .RN(rst_n), .Q(
        y_out_sum2[30]) );
  DFFRHQX1 y_out_sum6_reg_39_ ( .D(n3671), .CK(clk), .RN(rst_n), .Q(
        y_out_sum6[39]) );
  DFFRHQXL y_out_sum14_reg_29_ ( .D(n3201), .CK(clk), .RN(rst_n), .Q(
        y_out_sum14[29]) );
  DFFRHQX1 y_out_sum1_reg_19_ ( .D(n3917), .CK(clk), .RN(rst_n), .Q(
        y_out_sum1[19]) );
  DFFRHQX1 y_out_sum2_reg_15_ ( .D(n3875), .CK(clk), .RN(rst_n), .Q(
        y_out_sum2[15]) );
  DFFRHQXL y_out_sum2_reg_31_ ( .D(n3859), .CK(clk), .RN(rst_n), .Q(
        y_out_sum2[31]) );
  DFFRHQXL y_out_sum4_reg_33_ ( .D(n3747), .CK(clk), .RN(rst_n), .Q(
        y_out_sum4[33]) );
  DFFRHQX1 y_out_sum5_reg_13_ ( .D(n3712), .CK(clk), .RN(rst_n), .Q(
        y_out_sum5[13]) );
  DFFRHQX1 y_out_sum2_reg_16_ ( .D(n3874), .CK(clk), .RN(rst_n), .Q(
        y_out_sum2[16]) );
  DFFRHQX1 y_out_sum1_reg_16_ ( .D(n3920), .CK(clk), .RN(rst_n), .Q(
        y_out_sum1[16]) );
  DFFRHQX1 reg_length5_reg_5_ ( .D(n3672), .CK(clk), .RN(rst_n), .Q(
        reg_length5[5]) );
  DFFRX1 y_out_sum12_reg_14_ ( .D(n3326), .CK(clk), .RN(rst_n), .Q(
        y_out_sum12[14]), .QN(n4943) );
  DFFRHQX1 y_out_sum14_reg_16_ ( .D(n3214), .CK(clk), .RN(rst_n), .Q(
        y_out_sum14[16]) );
  DFFRHQX1 y_out_sum1_reg_18_ ( .D(n3918), .CK(clk), .RN(rst_n), .Q(
        y_out_sum1[18]) );
  DFFRHQXL y_out_sum4_reg_36_ ( .D(n3744), .CK(clk), .RN(rst_n), .Q(
        y_out_sum4[36]) );
  DFFRHQX1 y_out_sum2_reg_18_ ( .D(n3872), .CK(clk), .RN(rst_n), .Q(
        y_out_sum2[18]) );
  DFFRXL y_out_sum8_reg_27_ ( .D(n3533), .CK(clk), .RN(rst_n), .Q(
        y_out_sum8[27]), .QN(n6680) );
  DFFRHQXL y_out_sum11_reg_29_ ( .D(n3366), .CK(clk), .RN(rst_n), .Q(
        y_out_sum11[29]) );
  DFFRHQXL y_out_sum4_reg_32_ ( .D(n3748), .CK(clk), .RN(rst_n), .Q(
        y_out_sum4[32]) );
  DFFRHQXL y_out_sum5_reg_29_ ( .D(n3696), .CK(clk), .RN(rst_n), .Q(
        y_out_sum5[29]) );
  DFFRHQXL y_out_sum4_reg_37_ ( .D(n3743), .CK(clk), .RN(rst_n), .Q(
        y_out_sum4[37]) );
  DFFRHQX1 y_out_sum8_reg_12_ ( .D(n3548), .CK(clk), .RN(rst_n), .Q(
        y_out_sum8[12]) );
  DFFRHQX1 y_out_sum3_reg_12_ ( .D(n3823), .CK(clk), .RN(rst_n), .Q(
        y_out_sum3[12]) );
  DFFRHQX1 y_out_sum2_reg_21_ ( .D(n3869), .CK(clk), .RN(rst_n), .Q(
        y_out_sum2[21]) );
  DFFRHQXL y_out_sum2_reg_28_ ( .D(n3862), .CK(clk), .RN(rst_n), .Q(
        y_out_sum2[28]) );
  DFFRHQX1 y_out_sum11_reg_16_ ( .D(n3379), .CK(clk), .RN(rst_n), .Q(
        y_out_sum11[16]) );
  DFFRHQX1 y_out_sum2_reg_19_ ( .D(n3871), .CK(clk), .RN(rst_n), .Q(
        y_out_sum2[19]) );
  DFFRHQX1 y_out_sum2_reg_26_ ( .D(n3864), .CK(clk), .RN(rst_n), .Q(
        y_out_sum2[26]) );
  DFFRHQX1 y_out_sum4_reg_39_ ( .D(n3781), .CK(clk), .RN(rst_n), .Q(
        y_out_sum4[39]) );
  DFFRHQXL y_out_sum14_reg_28_ ( .D(n3202), .CK(clk), .RN(rst_n), .Q(
        y_out_sum14[28]) );
  DFFRHQX1 reg_length8_reg_4_ ( .D(n3508), .CK(clk), .RN(rst_n), .Q(
        reg_length8[4]) );
  DFFRX1 y_out_sum10_reg_14_ ( .D(n3436), .CK(clk), .RN(rst_n), .Q(
        y_out_sum10[14]), .QN(n4929) );
  DFFRX1 y_out_sum9_reg_14_ ( .D(n3491), .CK(clk), .RN(rst_n), .Q(
        y_out_sum9[14]), .QN(n4938) );
  DFFRHQX1 y_out_sum14_reg_21_ ( .D(n3209), .CK(clk), .RN(rst_n), .Q(
        y_out_sum14[21]) );
  DFFRHQX1 y_out_sum1_reg_20_ ( .D(n3916), .CK(clk), .RN(rst_n), .Q(
        y_out_sum1[20]) );
  DFFRHQXL y_out_sum5_reg_27_ ( .D(n3698), .CK(clk), .RN(rst_n), .Q(
        y_out_sum5[27]) );
  DFFRX1 y_out_sum12_reg_15_ ( .D(n3325), .CK(clk), .RN(rst_n), .Q(
        y_out_sum12[15]), .QN(n4891) );
  DFFRHQX1 y_out_sum5_reg_15_ ( .D(n3710), .CK(clk), .RN(rst_n), .Q(
        y_out_sum5[15]) );
  DFFRX1 y_out_sum13_reg_14_ ( .D(n3271), .CK(clk), .RN(rst_n), .Q(
        y_out_sum13[14]), .QN(n4940) );
  DFFRHQXL y_out_sum5_reg_31_ ( .D(n3694), .CK(clk), .RN(rst_n), .Q(
        y_out_sum5[31]) );
  DFFRHQXL y_out_sum11_reg_28_ ( .D(n3367), .CK(clk), .RN(rst_n), .Q(
        y_out_sum11[28]) );
  DFFRHQX1 reg_length2_reg_4_ ( .D(n3838), .CK(clk), .RN(rst_n), .Q(
        reg_length2[4]) );
  DFFRHQX1 y_out_sum11_reg_21_ ( .D(n3374), .CK(clk), .RN(rst_n), .Q(
        y_out_sum11[21]) );
  DFFRHQX1 y_out_sum10_reg_12_ ( .D(n3438), .CK(clk), .RN(rst_n), .Q(
        y_out_sum10[12]) );
  DFFRHQX1 y_out_sum7_reg_12_ ( .D(n3603), .CK(clk), .RN(rst_n), .Q(
        y_out_sum7[12]) );
  DFFRX1 y_out_sum7_reg_14_ ( .D(n3601), .CK(clk), .RN(rst_n), .Q(
        y_out_sum7[14]), .QN(n4931) );
  DFFRX1 y_out_sum9_reg_15_ ( .D(n3490), .CK(clk), .RN(rst_n), .Q(
        y_out_sum9[15]), .QN(n4885) );
  DFFRXL y_out_sum14_reg_30_ ( .D(n3200), .CK(clk), .RN(rst_n), .Q(
        y_out_sum14[30]), .QN(n6348) );
  DFFRX1 y_out_sum10_reg_15_ ( .D(n3435), .CK(clk), .RN(rst_n), .Q(
        y_out_sum10[15]), .QN(n4879) );
  DFFRHQX1 y_out_sum5_reg_12_ ( .D(n3713), .CK(clk), .RN(rst_n), .Q(
        y_out_sum5[12]) );
  DFFRHQX1 y_out_sum14_reg_20_ ( .D(n3210), .CK(clk), .RN(rst_n), .Q(
        y_out_sum14[20]) );
  DFFRHQX1 y_out_sum5_reg_14_ ( .D(n3711), .CK(clk), .RN(rst_n), .Q(
        y_out_sum5[14]) );
  DFFRHQX1 y_out_sum5_reg_17_ ( .D(n3708), .CK(clk), .RN(rst_n), .Q(
        y_out_sum5[17]) );
  DFFRHQX1 y_out_sum2_reg_12_ ( .D(n3878), .CK(clk), .RN(rst_n), .Q(
        y_out_sum2[12]) );
  DFFRX1 y_out_sum13_reg_15_ ( .D(n3270), .CK(clk), .RN(rst_n), .Q(
        y_out_sum13[15]), .QN(n4888) );
  DFFRHQXL y_out_sum5_reg_30_ ( .D(n3695), .CK(clk), .RN(rst_n), .Q(
        y_out_sum5[30]) );
  DFFRHQX1 y_out_sum2_reg_20_ ( .D(n3870), .CK(clk), .RN(rst_n), .Q(
        y_out_sum2[20]) );
  DFFRHQXL y_out_sum5_reg_28_ ( .D(n3697), .CK(clk), .RN(rst_n), .Q(
        y_out_sum5[28]) );
  DFFRHQX1 y_out_sum5_reg_21_ ( .D(n3704), .CK(clk), .RN(rst_n), .Q(
        y_out_sum5[21]) );
  DFFRHQX1 y_out_sum11_reg_20_ ( .D(n3375), .CK(clk), .RN(rst_n), .Q(
        y_out_sum11[20]) );
  DFFRX1 y_out_sum8_reg_18_ ( .D(n3542), .CK(clk), .RN(rst_n), .Q(
        y_out_sum8[18]), .QN(n4916) );
  DFFRHQX1 y_out_sum14_reg_13_ ( .D(n3217), .CK(clk), .RN(rst_n), .Q(
        y_out_sum14[13]) );
  DFFRXL y_out_sum11_reg_30_ ( .D(n3365), .CK(clk), .RN(rst_n), .Q(
        y_out_sum11[30]), .QN(n6509) );
  DFFRHQXL reg_length0_reg_5_ ( .D(n4028), .CK(clk), .RN(rst_n), .Q(
        reg_length0[5]) );
  DFFRHQX1 reg_length14_reg_5_ ( .D(n3177), .CK(clk), .RN(rst_n), .Q(
        reg_length14[5]) );
  DFFRX1 y_out_sum7_reg_15_ ( .D(n3600), .CK(clk), .RN(rst_n), .Q(
        y_out_sum7[15]), .QN(n4878) );
  DFFRHQX1 y_out_sum5_reg_11_ ( .D(n3714), .CK(clk), .RN(rst_n), .Q(
        y_out_sum5[11]) );
  DFFRX1 y_out_sum14_reg_22_ ( .D(n3208), .CK(clk), .RN(rst_n), .Q(
        y_out_sum14[22]), .QN(n4962) );
  DFFRHQX1 y_out_sum11_reg_13_ ( .D(n3382), .CK(clk), .RN(rst_n), .Q(
        y_out_sum11[13]) );
  DFFRHQX1 reg_length12_reg_3_ ( .D(n3289), .CK(clk), .RN(rst_n), .Q(
        reg_length12[3]) );
  DFFRXL y_out_sum14_reg_31_ ( .D(n3199), .CK(clk), .RN(rst_n), .Q(
        y_out_sum14[31]), .QN(n6346) );
  DFFRHQX1 y_out_sum13_reg_12_ ( .D(n3273), .CK(clk), .RN(rst_n), .Q(
        y_out_sum13[12]) );
  DFFRHQX1 y_out_sum5_reg_19_ ( .D(n3706), .CK(clk), .RN(rst_n), .Q(
        y_out_sum5[19]) );
  DFFRHQX1 reg_length1_reg_4_ ( .D(n3893), .CK(clk), .RN(rst_n), .Q(
        reg_length1[4]) );
  DFFRHQX1 y_out_sum6_reg_13_ ( .D(n3657), .CK(clk), .RN(rst_n), .Q(
        y_out_sum6[13]) );
  DFFRX1 y_out_sum8_reg_19_ ( .D(n3541), .CK(clk), .RN(rst_n), .Q(
        y_out_sum8[19]), .QN(n4865) );
  DFFRHQX1 y_out_sum0_reg_11_ ( .D(n3965), .CK(clk), .RN(rst_n), .Q(
        y_out_sum0[11]) );
  DFFRHQXL reg_length0_reg_4_ ( .D(n3990), .CK(clk), .RN(rst_n), .Q(
        reg_length0[4]) );
  DFFRHQX1 count_reg_7_ ( .D(n4019), .CK(clk), .RN(rst_n), .Q(N5060) );
  DFFRHQX1 reg_length6_reg_5_ ( .D(n3617), .CK(clk), .RN(rst_n), .Q(
        reg_length6[5]) );
  DFFRHQX1 reg_length9_reg_3_ ( .D(n3454), .CK(clk), .RN(rst_n), .Q(
        reg_length9[3]) );
  DFFRHQX1 y_out_sum5_reg_16_ ( .D(n3709), .CK(clk), .RN(rst_n), .Q(
        y_out_sum5[16]) );
  DFFRHQXL y_out_sum6_reg_29_ ( .D(n3641), .CK(clk), .RN(rst_n), .Q(
        y_out_sum6[29]) );
  DFFRXL y_out_sum11_reg_31_ ( .D(n3364), .CK(clk), .RN(rst_n), .Q(
        y_out_sum11[31]), .QN(n6507) );
  DFFRX1 y_out_sum11_reg_26_ ( .D(n3369), .CK(clk), .RN(rst_n), .Q(
        y_out_sum11[26]), .QN(n4960) );
  DFFRHQX1 y_out_sum5_reg_18_ ( .D(n3707), .CK(clk), .RN(rst_n), .Q(
        y_out_sum5[18]) );
  DFFRHQX1 y_out_sum1_reg_12_ ( .D(n3924), .CK(clk), .RN(rst_n), .Q(
        y_out_sum1[12]) );
  DFFRHQX1 y_out_sum12_reg_12_ ( .D(n3328), .CK(clk), .RN(rst_n), .Q(
        y_out_sum12[12]) );
  DFFRXL y_out_sum14_reg_27_ ( .D(n3203), .CK(clk), .RN(rst_n), .Q(
        y_out_sum14[27]), .QN(n6352) );
  DFFRHQX1 y_out_sum14_reg_12_ ( .D(n3218), .CK(clk), .RN(rst_n), .Q(
        y_out_sum14[12]) );
  DFFRHQX1 y_out_sum4_reg_13_ ( .D(n3767), .CK(clk), .RN(rst_n), .Q(
        y_out_sum4[13]) );
  DFFRHQX1 reg_length11_reg_5_ ( .D(n3342), .CK(clk), .RN(rst_n), .Q(
        reg_length11[5]) );
  DFFRHQX1 y_out_sum5_reg_20_ ( .D(n3705), .CK(clk), .RN(rst_n), .Q(
        y_out_sum5[20]) );
  DFFRHQX1 y_out_sum6_reg_15_ ( .D(n3655), .CK(clk), .RN(rst_n), .Q(
        y_out_sum6[15]) );
  DFFRHQXL y_out_sum6_reg_31_ ( .D(n3639), .CK(clk), .RN(rst_n), .Q(
        y_out_sum6[31]) );
  DFFRHQX1 reg_length4_reg_5_ ( .D(n3727), .CK(clk), .RN(rst_n), .Q(
        reg_length4[5]) );
  DFFRX1 y_out_sum14_reg_23_ ( .D(n3207), .CK(clk), .RN(rst_n), .Q(
        y_out_sum14[23]), .QN(n4957) );
  DFFRHQXL y_out_sum6_reg_27_ ( .D(n3643), .CK(clk), .RN(rst_n), .Q(
        y_out_sum6[27]) );
  DFFRXL y_out_sum11_reg_27_ ( .D(n3368), .CK(clk), .RN(rst_n), .Q(
        y_out_sum11[27]), .QN(n6513) );
  DFFRHQXL y_out_sum4_reg_29_ ( .D(n3751), .CK(clk), .RN(rst_n), .Q(
        y_out_sum4[29]) );
  DFFRHQX1 y_out_sum11_reg_12_ ( .D(n3383), .CK(clk), .RN(rst_n), .Q(
        y_out_sum11[12]) );
  DFFRHQX1 reg_length13_reg_3_ ( .D(n3234), .CK(clk), .RN(rst_n), .Q(
        reg_length13[3]) );
  DFFRHQX1 reg_length5_reg_4_ ( .D(n3673), .CK(clk), .RN(rst_n), .Q(
        reg_length5[4]) );
  DFFRHQX1 reg_length14_reg_4_ ( .D(n3178), .CK(clk), .RN(rst_n), .Q(
        reg_length14[4]) );
  DFFRHQX1 y_out_sum6_reg_14_ ( .D(n3656), .CK(clk), .RN(rst_n), .Q(
        y_out_sum6[14]) );
  DFFRHQX1 y_out_sum6_reg_12_ ( .D(n3658), .CK(clk), .RN(rst_n), .Q(
        y_out_sum6[12]) );
  DFFRHQXL y_out_sum4_reg_27_ ( .D(n3753), .CK(clk), .RN(rst_n), .Q(
        y_out_sum4[27]) );
  DFFRHQX1 reg_length7_reg_3_ ( .D(n3564), .CK(clk), .RN(rst_n), .Q(
        reg_length7[3]) );
  DFFRHQX1 y_out_sum6_reg_17_ ( .D(n3653), .CK(clk), .RN(rst_n), .Q(
        y_out_sum6[17]) );
  DFFRHQX1 y_out_sum4_reg_15_ ( .D(n3765), .CK(clk), .RN(rst_n), .Q(
        y_out_sum4[15]) );
  DFFRHQX1 y_out_sum3_reg_11_ ( .D(n3824), .CK(clk), .RN(rst_n), .Q(
        y_out_sum3[11]) );
  DFFRHQX1 reg_length11_reg_4_ ( .D(n3343), .CK(clk), .RN(rst_n), .Q(
        reg_length11[4]) );
  DFFRHQXL y_out_sum6_reg_30_ ( .D(n3640), .CK(clk), .RN(rst_n), .Q(
        y_out_sum6[30]) );
  DFFRHQXL y_out_sum4_reg_31_ ( .D(n3749), .CK(clk), .RN(rst_n), .Q(
        y_out_sum4[31]) );
  DFFRHQX1 y_out_sum2_reg_11_ ( .D(n3879), .CK(clk), .RN(rst_n), .Q(
        y_out_sum2[11]) );
  DFFRHQXL y_out_sum6_reg_28_ ( .D(n3642), .CK(clk), .RN(rst_n), .Q(
        y_out_sum6[28]) );
  DFFRHQX1 y_out_sum6_reg_21_ ( .D(n3649), .CK(clk), .RN(rst_n), .Q(
        y_out_sum6[21]) );
  DFFRHQX1 y_out_sum4_reg_14_ ( .D(n3766), .CK(clk), .RN(rst_n), .Q(
        y_out_sum4[14]) );
  DFFRX1 y_out_sum8_reg_14_ ( .D(n3546), .CK(clk), .RN(rst_n), .Q(
        y_out_sum8[14]), .QN(n4919) );
  DFFRHQX1 y_out_sum4_reg_11_ ( .D(n3769), .CK(clk), .RN(rst_n), .Q(
        y_out_sum4[11]) );
  DFFRHQX1 y_out_sum6_reg_26_ ( .D(n3644), .CK(clk), .RN(rst_n), .Q(
        y_out_sum6[26]) );
  DFFRHQX1 y_out_sum4_reg_12_ ( .D(n3768), .CK(clk), .RN(rst_n), .Q(
        y_out_sum4[12]) );
  DFFRX1 y_out_sum14_reg_18_ ( .D(n3212), .CK(clk), .RN(rst_n), .Q(
        y_out_sum14[18]), .QN(n4910) );
  DFFRHQX1 y_out_sum6_reg_19_ ( .D(n3651), .CK(clk), .RN(rst_n), .Q(
        y_out_sum6[19]) );
  DFFRHQX1 y_out_sum4_reg_17_ ( .D(n3763), .CK(clk), .RN(rst_n), .Q(
        y_out_sum4[17]) );
  DFFRHQXL y_out_sum4_reg_30_ ( .D(n3750), .CK(clk), .RN(rst_n), .Q(
        y_out_sum4[30]) );
  DFFRHQX1 y_out_sum5_reg_10_ ( .D(n3715), .CK(clk), .RN(rst_n), .Q(
        y_out_sum5[10]) );
  DFFRHQX1 y_out_sum6_reg_11_ ( .D(n3659), .CK(clk), .RN(rst_n), .Q(
        y_out_sum6[11]) );
  DFFRHQXL y_out_sum4_reg_28_ ( .D(n3752), .CK(clk), .RN(rst_n), .Q(
        y_out_sum4[28]) );
  DFFRHQX1 y_out_sum6_reg_16_ ( .D(n3654), .CK(clk), .RN(rst_n), .Q(
        y_out_sum6[16]) );
  DFFRHQX1 y_out_sum4_reg_21_ ( .D(n3759), .CK(clk), .RN(rst_n), .Q(
        y_out_sum4[21]) );
  DFFRX1 y_out_sum11_reg_18_ ( .D(n3377), .CK(clk), .RN(rst_n), .Q(
        y_out_sum11[18]), .QN(n4905) );
  DFFRX1 y_out_sum8_reg_15_ ( .D(n3545), .CK(clk), .RN(rst_n), .Q(
        y_out_sum8[15]), .QN(n4866) );
  DFFRHQX1 reg_length10_reg_3_ ( .D(n3399), .CK(clk), .RN(rst_n), .Q(
        reg_length10[3]) );
  DFFRHQX1 y_out_sum6_reg_18_ ( .D(n3652), .CK(clk), .RN(rst_n), .Q(
        y_out_sum6[18]) );
  DFFRX1 y_out_sum14_reg_19_ ( .D(n3211), .CK(clk), .RN(rst_n), .Q(
        y_out_sum14[19]), .QN(n4859) );
  DFFRHQX1 y_out_sum4_reg_19_ ( .D(n3761), .CK(clk), .RN(rst_n), .Q(
        y_out_sum4[19]) );
  DFFRX1 y_out_sum11_reg_19_ ( .D(n3376), .CK(clk), .RN(rst_n), .Q(
        y_out_sum11[19]), .QN(n4854) );
  DFFRHQX1 y_out_sum6_reg_20_ ( .D(n3650), .CK(clk), .RN(rst_n), .Q(
        y_out_sum6[20]) );
  DFFRHQX1 y_out_sum4_reg_16_ ( .D(n3764), .CK(clk), .RN(rst_n), .Q(
        y_out_sum4[16]) );
  DFFRHQX1 y_out_sum1_reg_11_ ( .D(n3925), .CK(clk), .RN(rst_n), .Q(
        y_out_sum1[11]) );
  DFFRX1 y_out_sum8_reg_11_ ( .D(n3549), .CK(clk), .RN(rst_n), .Q(
        y_out_sum8[11]), .QN(n4864) );
  DFFRHQX1 y_out_sum4_reg_18_ ( .D(n3762), .CK(clk), .RN(rst_n), .Q(
        y_out_sum4[18]) );
  DFFRHQX1 y_out_sum0_reg_10_ ( .D(n3966), .CK(clk), .RN(rst_n), .Q(
        y_out_sum0[10]) );
  DFFRX1 y_out_sum10_reg_11_ ( .D(n3439), .CK(clk), .RN(rst_n), .Q(
        y_out_sum10[11]), .QN(n4876) );
  DFFRX1 y_out_sum9_reg_11_ ( .D(n3494), .CK(clk), .RN(rst_n), .Q(
        y_out_sum9[11]), .QN(n4881) );
  DFFRHQX1 y_out_sum4_reg_20_ ( .D(n3760), .CK(clk), .RN(rst_n), .Q(
        y_out_sum4[20]) );
  DFFRX1 y_out_sum7_reg_11_ ( .D(n3604), .CK(clk), .RN(rst_n), .Q(
        y_out_sum7[11]), .QN(n4875) );
  DFFRHQX1 y_out_sum3_reg_10_ ( .D(n3825), .CK(clk), .RN(rst_n), .Q(
        y_out_sum3[10]) );
  DFFRHQXL reg_length0_reg_3_ ( .D(n3989), .CK(clk), .RN(rst_n), .Q(
        reg_length0[3]) );
  DFFRHQX1 y_out_sum4_reg_10_ ( .D(n3770), .CK(clk), .RN(rst_n), .Q(
        y_out_sum4[10]) );
  DFFRHQX1 y_out_sum2_reg_10_ ( .D(n3880), .CK(clk), .RN(rst_n), .Q(
        y_out_sum2[10]) );
  DFFRHQX1 reg_length8_reg_3_ ( .D(n3509), .CK(clk), .RN(rst_n), .Q(
        reg_length8[3]) );
  DFFRHQX1 reg_length9_reg_2_ ( .D(n3455), .CK(clk), .RN(rst_n), .Q(
        reg_length9[2]) );
  DFFRX1 y_out_sum14_reg_14_ ( .D(n3216), .CK(clk), .RN(rst_n), .Q(
        y_out_sum14[14]), .QN(n4912) );
  DFFRHQX1 reg_length6_reg_4_ ( .D(n3618), .CK(clk), .RN(rst_n), .Q(
        reg_length6[4]) );
  DFFRHQX1 y_out_sum6_reg_10_ ( .D(n3660), .CK(clk), .RN(rst_n), .Q(
        y_out_sum6[10]) );
  DFFRX1 y_out_sum11_reg_14_ ( .D(n3381), .CK(clk), .RN(rst_n), .Q(
        y_out_sum11[14]), .QN(n4909) );
  DFFRX1 y_out_sum12_reg_11_ ( .D(n3329), .CK(clk), .RN(rst_n), .Q(
        y_out_sum12[11]), .QN(n4890) );
  DFFRX1 y_out_sum8_reg_10_ ( .D(n3550), .CK(clk), .RN(rst_n), .Q(
        y_out_sum8[10]), .QN(n4915) );
  DFFRX1 y_out_sum13_reg_11_ ( .D(n3274), .CK(clk), .RN(rst_n), .Q(
        y_out_sum13[11]), .QN(n4886) );
  DFFRX1 y_out_sum14_reg_15_ ( .D(n3215), .CK(clk), .RN(rst_n), .Q(
        y_out_sum14[15]), .QN(n4861) );
  DFFRHQX1 reg_length4_reg_4_ ( .D(n3728), .CK(clk), .RN(rst_n), .Q(
        reg_length4[4]) );
  DFFRX1 y_out_sum11_reg_15_ ( .D(n3380), .CK(clk), .RN(rst_n), .Q(
        y_out_sum11[15]), .QN(n4857) );
  DFFRX1 y_out_sum14_reg_11_ ( .D(n3219), .CK(clk), .RN(rst_n), .Q(
        y_out_sum14[11]), .QN(n4860) );
  DFFRHQX1 y_out_sum1_reg_10_ ( .D(n3926), .CK(clk), .RN(rst_n), .Q(
        y_out_sum1[10]) );
  DFFRX1 y_out_sum11_reg_11_ ( .D(n3384), .CK(clk), .RN(rst_n), .Q(
        y_out_sum11[11]), .QN(n4856) );
  DFFRHQX1 reg_length13_reg_2_ ( .D(n3235), .CK(clk), .RN(rst_n), .Q(
        reg_length13[2]) );
  DFFRX1 y_out_sum10_reg_10_ ( .D(n3440), .CK(clk), .RN(rst_n), .Q(
        y_out_sum10[10]), .QN(n4928) );
  DFFRHQX1 reg_length12_reg_2_ ( .D(n3290), .CK(clk), .RN(rst_n), .Q(
        reg_length12[2]) );
  DFFRHQX1 reg_length10_reg_2_ ( .D(n3400), .CK(clk), .RN(rst_n), .Q(
        reg_length10[2]) );
  DFFRHQX1 y_out_sum5_reg_9_ ( .D(n3716), .CK(clk), .RN(rst_n), .Q(
        y_out_sum5[9]) );
  DFFRHQX1 reg_length14_reg_3_ ( .D(n3179), .CK(clk), .RN(rst_n), .Q(
        reg_length14[3]) );
  DFFRX1 y_out_sum7_reg_10_ ( .D(n3605), .CK(clk), .RN(rst_n), .Q(
        y_out_sum7[10]), .QN(n4926) );
  DFFRHQX1 y_out_sum8_reg_9_ ( .D(n3551), .CK(clk), .RN(rst_n), .Q(
        y_out_sum8[9]) );
  DFFRHQX1 y_out_sum0_reg_9_ ( .D(n3967), .CK(clk), .RN(rst_n), .Q(
        y_out_sum0[9]) );
  DFFRX1 y_out_sum13_reg_10_ ( .D(n3275), .CK(clk), .RN(rst_n), .Q(
        y_out_sum13[10]), .QN(n4939) );
  DFFRHQX1 reg_length7_reg_2_ ( .D(n3565), .CK(clk), .RN(rst_n), .Q(
        reg_length7[2]) );
  DFFRX1 y_out_sum14_reg_10_ ( .D(n3220), .CK(clk), .RN(rst_n), .Q(
        y_out_sum14[10]), .QN(n4911) );
  DFFRX1 y_out_sum9_reg_10_ ( .D(n3495), .CK(clk), .RN(rst_n), .Q(
        y_out_sum9[10]), .QN(n4932) );
  DFFRHQX1 reg_length11_reg_3_ ( .D(n3344), .CK(clk), .RN(rst_n), .Q(
        reg_length11[3]) );
  DFFRX1 y_out_sum12_reg_10_ ( .D(n3330), .CK(clk), .RN(rst_n), .Q(
        y_out_sum12[10]), .QN(n4942) );
  DFFRX1 y_out_sum11_reg_10_ ( .D(n3385), .CK(clk), .RN(rst_n), .Q(
        y_out_sum11[10]), .QN(n4908) );
  DFFRHQX1 y_out_sum2_reg_9_ ( .D(n3881), .CK(clk), .RN(rst_n), .Q(
        y_out_sum2[9]) );
  DFFRHQX1 y_out_sum9_reg_9_ ( .D(n3496), .CK(clk), .RN(rst_n), .Q(
        y_out_sum9[9]) );
  DFFRHQX1 count_reg_4_ ( .D(n4022), .CK(clk), .RN(rst_n), .Q(count[4]) );
  DFFRHQX1 y_out_sum4_reg_9_ ( .D(n3771), .CK(clk), .RN(rst_n), .Q(
        y_out_sum4[9]) );
  DFFRHQX1 y_out_sum7_reg_9_ ( .D(n3606), .CK(clk), .RN(rst_n), .Q(
        y_out_sum7[9]) );
  DFFRHQX1 y_out_sum14_reg_9_ ( .D(n3221), .CK(clk), .RN(rst_n), .Q(
        y_out_sum14[9]) );
  DFFRHQX1 count_reg_6_ ( .D(n4020), .CK(clk), .RN(rst_n), .Q(N5059) );
  DFFRHQX1 y_out_sum13_reg_9_ ( .D(n3276), .CK(clk), .RN(rst_n), .Q(
        y_out_sum13[9]) );
  DFFRHQX1 y_out_sum10_reg_9_ ( .D(n3441), .CK(clk), .RN(rst_n), .Q(
        y_out_sum10[9]) );
  DFFRHQX1 reg_length8_reg_2_ ( .D(n3510), .CK(clk), .RN(rst_n), .Q(
        reg_length8[2]) );
  DFFRHQX1 count_reg_5_ ( .D(n4021), .CK(clk), .RN(rst_n), .Q(N5058) );
  DFFRHQX1 y_out_sum0_reg_8_ ( .D(n3968), .CK(clk), .RN(rst_n), .Q(
        y_out_sum0[8]) );
  DFFRHQX1 y_out_sum11_reg_9_ ( .D(n3386), .CK(clk), .RN(rst_n), .Q(
        y_out_sum11[9]) );
  DFFRHQX1 y_out_sum8_reg_8_ ( .D(n3552), .CK(clk), .RN(rst_n), .Q(
        y_out_sum8[8]) );
  DFFRHQX1 y_out_sum1_reg_9_ ( .D(n3927), .CK(clk), .RN(rst_n), .Q(
        y_out_sum1[9]) );
  DFFRHQX1 count_reg_3_ ( .D(n4023), .CK(clk), .RN(rst_n), .Q(count[3]) );
  DFFRHQX1 y_out_sum12_reg_9_ ( .D(n3331), .CK(clk), .RN(rst_n), .Q(
        y_out_sum12[9]) );
  DFFRHQX1 y_out_sum3_reg_9_ ( .D(n3826), .CK(clk), .RN(rst_n), .Q(
        y_out_sum3[9]) );
  DFFRHQX1 y_out_sum5_reg_8_ ( .D(n3717), .CK(clk), .RN(rst_n), .Q(
        y_out_sum5[8]) );
  DFFRHQX1 reg_length0_reg_0_ ( .D(n3991), .CK(clk), .RN(rst_n), .Q(
        reg_length0[0]) );
  DFFRHQX1 y_out_sum6_reg_9_ ( .D(n3661), .CK(clk), .RN(rst_n), .Q(
        y_out_sum6[9]) );
  DFFRHQX1 count_reg_2_ ( .D(n4024), .CK(clk), .RN(rst_n), .Q(count[2]) );
  DFFRHQX1 y_out_sum13_reg_8_ ( .D(n3277), .CK(clk), .RN(rst_n), .Q(
        y_out_sum13[8]) );
  DFFRHQX1 y_out_sum2_reg_8_ ( .D(n3882), .CK(clk), .RN(rst_n), .Q(
        y_out_sum2[8]) );
  DFFRHQX1 count_reg_0_ ( .D(n4025), .CK(clk), .RN(rst_n), .Q(count[0]) );
  DFFRHQX1 reg_length14_reg_2_ ( .D(n3180), .CK(clk), .RN(rst_n), .Q(
        reg_length14[2]) );
  DFFRHQX1 y_out_sum4_reg_8_ ( .D(n3772), .CK(clk), .RN(rst_n), .Q(
        y_out_sum4[8]) );
  DFFRHQX1 y_out_sum3_reg_8_ ( .D(n3827), .CK(clk), .RN(rst_n), .Q(
        y_out_sum3[8]) );
  DFFRHQX1 y_out_sum14_reg_8_ ( .D(n3222), .CK(clk), .RN(rst_n), .Q(
        y_out_sum14[8]) );
  DFFRHQX1 count_reg_1_ ( .D(n4026), .CK(clk), .RN(rst_n), .Q(count[1]) );
  DFFRHQX1 y_out_sum7_reg_8_ ( .D(n3607), .CK(clk), .RN(rst_n), .Q(
        y_out_sum7[8]) );
  DFFRHQX1 reg_length11_reg_2_ ( .D(n3345), .CK(clk), .RN(rst_n), .Q(
        reg_length11[2]) );
  DFFRHQX1 y_out_sum12_reg_8_ ( .D(n3332), .CK(clk), .RN(rst_n), .Q(
        y_out_sum12[8]) );
  DFFRHQX1 reg_length3_reg_3_ ( .D(n3784), .CK(clk), .RN(rst_n), .Q(
        reg_length3[3]) );
  DFFRHQX1 reg_length9_reg_1_ ( .D(n3456), .CK(clk), .RN(rst_n), .Q(
        reg_length9[1]) );
  DFFRHQX1 y_out_sum6_reg_8_ ( .D(n3662), .CK(clk), .RN(rst_n), .Q(
        y_out_sum6[8]) );
  DFFRHQX1 y_out_sum9_reg_8_ ( .D(n3497), .CK(clk), .RN(rst_n), .Q(
        y_out_sum9[8]) );
  DFFRHQX1 y_out_sum10_reg_8_ ( .D(n3442), .CK(clk), .RN(rst_n), .Q(
        y_out_sum10[8]) );
  DFFRHQX1 y_out_sum0_reg_7_ ( .D(n3969), .CK(clk), .RN(rst_n), .Q(
        y_out_sum0[7]) );
  DFFRHQX1 y_out_sum5_reg_7_ ( .D(n3718), .CK(clk), .RN(rst_n), .Q(
        y_out_sum5[7]) );
  DFFRHQX1 y_out_sum11_reg_8_ ( .D(n3387), .CK(clk), .RN(rst_n), .Q(
        y_out_sum11[8]) );
  DFFRHQX1 reg_length10_reg_1_ ( .D(n3401), .CK(clk), .RN(rst_n), .Q(
        reg_length10[1]) );
  DFFRHQX1 y_out_sum2_reg_7_ ( .D(n3883), .CK(clk), .RN(rst_n), .Q(
        y_out_sum2[7]) );
  DFFRHQX1 y_out_sum1_reg_8_ ( .D(n3928), .CK(clk), .RN(rst_n), .Q(
        y_out_sum1[8]) );
  DFFRHQX1 y_out_sum4_reg_7_ ( .D(n3773), .CK(clk), .RN(rst_n), .Q(
        y_out_sum4[7]) );
  DFFRHQX1 reg_length12_reg_1_ ( .D(n3291), .CK(clk), .RN(rst_n), .Q(
        reg_length12[1]) );
  DFFRHQX1 reg_length2_reg_3_ ( .D(n3839), .CK(clk), .RN(rst_n), .Q(
        reg_length2[3]) );
  DFFRHQX1 y_out_sum3_reg_7_ ( .D(n3828), .CK(clk), .RN(rst_n), .Q(
        y_out_sum3[7]) );
  DFFRHQX1 y_out_sum6_reg_7_ ( .D(n3663), .CK(clk), .RN(rst_n), .Q(
        y_out_sum6[7]) );
  DFFRHQX1 reg_length12_reg_0_ ( .D(n3292), .CK(clk), .RN(rst_n), .Q(
        reg_length12[0]) );
  DFFRHQX1 reg_length1_reg_3_ ( .D(n3894), .CK(clk), .RN(rst_n), .Q(
        reg_length1[3]) );
  DFFRX1 y_out_sum8_reg_7_ ( .D(n3553), .CK(clk), .RN(rst_n), .Q(y_out_sum8[7]), .QN(n4862) );
  DFFRHQX1 y_out_sum5_reg_6_ ( .D(n3719), .CK(clk), .RN(rst_n), .Q(
        y_out_sum5[6]) );
  DFFRHQX1 reg_length10_reg_0_ ( .D(n3402), .CK(clk), .RN(rst_n), .Q(
        reg_length10[0]) );
  DFFRHQX1 reg_length7_reg_1_ ( .D(n3566), .CK(clk), .RN(rst_n), .Q(
        reg_length7[1]) );
  DFFRHQX1 y_out_sum3_reg_6_ ( .D(n3829), .CK(clk), .RN(rst_n), .Q(
        y_out_sum3[6]) );
  DFFRHQX1 y_out_sum0_reg_6_ ( .D(n3970), .CK(clk), .RN(rst_n), .Q(
        y_out_sum0[6]) );
  DFFRHQX1 y_out_sum1_reg_7_ ( .D(n3929), .CK(clk), .RN(rst_n), .Q(
        y_out_sum1[7]) );
  DFFRHQX1 reg_length13_reg_0_ ( .D(n3237), .CK(clk), .RN(rst_n), .Q(
        reg_length13[0]) );
  DFFRHQX1 y_out_sum2_reg_6_ ( .D(n3884), .CK(clk), .RN(rst_n), .Q(
        y_out_sum2[6]) );
  DFFRHQX1 reg_length7_reg_0_ ( .D(n3567), .CK(clk), .RN(rst_n), .Q(
        reg_length7[0]) );
  DFFRHQX1 reg_length9_reg_0_ ( .D(n3457), .CK(clk), .RN(rst_n), .Q(
        reg_length9[0]) );
  DFFRHQX1 y_out_sum4_reg_6_ ( .D(n3774), .CK(clk), .RN(rst_n), .Q(
        y_out_sum4[6]) );
  DFFRX1 y_out_sum14_reg_7_ ( .D(n3223), .CK(clk), .RN(rst_n), .Q(
        y_out_sum14[7]), .QN(n4855) );
  DFFRX1 y_out_sum13_reg_7_ ( .D(n3278), .CK(clk), .RN(rst_n), .Q(
        y_out_sum13[7]), .QN(n4874) );
  DFFRHQX1 reg_length5_reg_3_ ( .D(n3674), .CK(clk), .RN(rst_n), .Q(
        reg_length5[3]) );
  DFFRX1 y_out_sum9_reg_7_ ( .D(n3498), .CK(clk), .RN(rst_n), .Q(y_out_sum9[7]), .QN(n4871) );
  DFFRHQX1 reg_length3_reg_2_ ( .D(n3785), .CK(clk), .RN(rst_n), .Q(
        reg_length3[2]) );
  DFFRX1 y_out_sum11_reg_7_ ( .D(n3388), .CK(clk), .RN(rst_n), .Q(
        y_out_sum11[7]), .QN(n4852) );
  DFFRHQX1 y_out_sum6_reg_6_ ( .D(n3664), .CK(clk), .RN(rst_n), .Q(
        y_out_sum6[6]) );
  DFFRX1 y_out_sum8_reg_6_ ( .D(n3554), .CK(clk), .RN(rst_n), .Q(y_out_sum8[6]), .QN(n4914) );
  DFFRHQX1 y_out_sum1_reg_6_ ( .D(n3930), .CK(clk), .RN(rst_n), .Q(
        y_out_sum1[6]) );
  DFFRX1 y_out_sum12_reg_7_ ( .D(n3333), .CK(clk), .RN(rst_n), .Q(
        y_out_sum12[7]), .QN(n4883) );
  DFFRHQX1 reg_length8_reg_1_ ( .D(n3511), .CK(clk), .RN(rst_n), .Q(
        reg_length8[1]) );
  DFFRX1 reg_length13_reg_1_ ( .D(n3236), .CK(clk), .RN(rst_n), .Q(
        reg_length13[1]), .QN(n4901) );
  DFFRHQX1 next_reg_0_ ( .D(n4009), .CK(clk), .RN(rst_n), .Q(next[0]) );
  DFFRX1 y_out_sum10_reg_7_ ( .D(n3443), .CK(clk), .RN(rst_n), .Q(
        y_out_sum10[7]), .QN(n4868) );
  DFFRX1 y_out_sum7_reg_7_ ( .D(n3608), .CK(clk), .RN(rst_n), .Q(y_out_sum7[7]), .QN(n4867) );
  DFFRHQX1 reg_length2_reg_2_ ( .D(n3840), .CK(clk), .RN(rst_n), .Q(
        reg_length2[2]) );
  DFFRX1 y_out_sum14_reg_6_ ( .D(n3224), .CK(clk), .RN(rst_n), .Q(
        y_out_sum14[6]), .QN(n4907) );
  DFFRX1 y_out_sum9_reg_6_ ( .D(n3499), .CK(clk), .RN(rst_n), .Q(y_out_sum9[6]), .QN(n4923) );
  DFFRHQX1 y_out_sum8_reg_5_ ( .D(n3555), .CK(clk), .RN(rst_n), .Q(
        y_out_sum8[5]) );
  DFFRHQX1 reg_length1_reg_2_ ( .D(n3895), .CK(clk), .RN(rst_n), .Q(
        reg_length1[2]) );
  DFFRHQX1 y_out_sum5_reg_5_ ( .D(n3720), .CK(clk), .RN(rst_n), .Q(
        y_out_sum5[5]) );
  DFFRHQX1 next_reg_1_ ( .D(n4027), .CK(clk), .RN(rst_n), .Q(next[1]) );
  DFFRHQX1 reg_length6_reg_3_ ( .D(n3619), .CK(clk), .RN(rst_n), .Q(
        reg_length6[3]) );
  DFFRX1 y_out_sum12_reg_6_ ( .D(n3334), .CK(clk), .RN(rst_n), .Q(
        y_out_sum12[6]), .QN(n4937) );
  DFFRHQX1 y_out_sum14_reg_5_ ( .D(n3225), .CK(clk), .RN(rst_n), .Q(
        y_out_sum14[5]) );
  DFFRX1 y_out_sum11_reg_6_ ( .D(n3389), .CK(clk), .RN(rst_n), .Q(
        y_out_sum11[6]), .QN(n4904) );
  DFFRHQX1 y_out_sum0_reg_5_ ( .D(n3971), .CK(clk), .RN(rst_n), .Q(
        y_out_sum0[5]) );
  DFFRHQX1 y_out_sum9_reg_5_ ( .D(n3500), .CK(clk), .RN(rst_n), .Q(
        y_out_sum9[5]) );
  DFFRX1 y_out_sum7_reg_6_ ( .D(n3609), .CK(clk), .RN(rst_n), .Q(y_out_sum7[6]), .QN(n4917) );
  DFFRX1 y_out_sum10_reg_6_ ( .D(n3444), .CK(clk), .RN(rst_n), .Q(
        y_out_sum10[6]), .QN(n4921) );
  DFFRHQXL out_value_reg ( .D(n2859), .CK(clk), .RN(rst_n), .Q(out_value) );
  DFFRHQX1 reg_length14_reg_1_ ( .D(n3181), .CK(clk), .RN(rst_n), .Q(
        reg_length14[1]) );
  DFFRHQX1 reg_length11_reg_1_ ( .D(n3346), .CK(clk), .RN(rst_n), .Q(
        reg_length11[1]) );
  DFFRHQX1 y_out_sum4_reg_5_ ( .D(n3775), .CK(clk), .RN(rst_n), .Q(
        y_out_sum4[5]) );
  DFFRHQX1 y_out_sum3_reg_5_ ( .D(n3830), .CK(clk), .RN(rst_n), .Q(
        y_out_sum3[5]) );
  DFFRHQX1 reg_length4_reg_3_ ( .D(n3729), .CK(clk), .RN(rst_n), .Q(
        reg_length4[3]) );
  DFFRX1 y_out_sum13_reg_6_ ( .D(n3279), .CK(clk), .RN(rst_n), .Q(
        y_out_sum13[6]), .QN(n4930) );
  DFFRHQX1 out_valid_reg ( .D(n3978), .CK(clk), .RN(rst_n), .Q(out_valid) );
  DFFRHQX1 reg_length3_reg_0_ ( .D(n3787), .CK(clk), .RN(rst_n), .Q(
        reg_length3[0]) );
  DFFRHQX1 reg_length5_reg_2_ ( .D(n3675), .CK(clk), .RN(rst_n), .Q(
        reg_length5[2]) );
  DFFRHQX1 reg_length3_reg_1_ ( .D(n3786), .CK(clk), .RN(rst_n), .Q(
        reg_length3[1]) );
  DFFRHQX1 y_out_sum2_reg_5_ ( .D(n3885), .CK(clk), .RN(rst_n), .Q(
        y_out_sum2[5]) );
  DFFRHQX1 y_out_sum11_reg_5_ ( .D(n3390), .CK(clk), .RN(rst_n), .Q(
        y_out_sum11[5]) );
  DFFRHQX1 y_out_sum12_reg_5_ ( .D(n3335), .CK(clk), .RN(rst_n), .Q(
        y_out_sum12[5]) );
  DFFRX1 next_reg_3_ ( .D(n4007), .CK(clk), .RN(rst_n), .Q(next[3]), .QN(n4849) );
  DFFRHQX1 y_out_sum6_reg_5_ ( .D(n3665), .CK(clk), .RN(rst_n), .Q(
        y_out_sum6[5]) );
  DFFRHQX1 y_out_sum10_reg_5_ ( .D(n3445), .CK(clk), .RN(rst_n), .Q(
        y_out_sum10[5]) );
  DFFRX1 reg_length8_reg_0_ ( .D(n3512), .CK(clk), .RN(rst_n), .Q(
        reg_length8[0]), .QN(n4902) );
  DFFRHQX1 y_out_sum13_reg_5_ ( .D(n3280), .CK(clk), .RN(rst_n), .Q(
        y_out_sum13[5]) );
  DFFRHQX1 reg_length11_reg_0_ ( .D(n3347), .CK(clk), .RN(rst_n), .Q(
        reg_length11[0]) );
  DFFRHQX1 y_out_sum7_reg_5_ ( .D(n3610), .CK(clk), .RN(rst_n), .Q(
        y_out_sum7[5]) );
  DFFRHQX1 y_out_sum1_reg_5_ ( .D(n3931), .CK(clk), .RN(rst_n), .Q(
        y_out_sum1[5]) );
  DFFRHQX1 reg_length2_reg_1_ ( .D(n3841), .CK(clk), .RN(rst_n), .Q(
        reg_length2[1]) );
  DFFRHQX1 reg_length1_reg_0_ ( .D(n3897), .CK(clk), .RN(rst_n), .Q(
        reg_length1[0]) );
  DFFRHQX1 reg_length1_reg_1_ ( .D(n3896), .CK(clk), .RN(rst_n), .Q(
        reg_length1[1]) );
  DFFRHQX1 y_out_sum5_reg_4_ ( .D(n3721), .CK(clk), .RN(rst_n), .Q(
        y_out_sum5[4]) );
  DFFRHQX1 next_reg_4_ ( .D(n4006), .CK(clk), .RN(rst_n), .Q(next[4]) );
  DFFRHQX1 next_reg_2_ ( .D(n4008), .CK(clk), .RN(rst_n), .Q(next[2]) );
  DFFRHQX1 y_out_sum3_reg_4_ ( .D(n3831), .CK(clk), .RN(rst_n), .Q(
        y_out_sum3[4]) );
  DFFRHQX1 reg_length2_reg_0_ ( .D(n3842), .CK(clk), .RN(rst_n), .Q(
        reg_length2[0]) );
  DFFRHQX1 y_out_sum0_reg_4_ ( .D(n3972), .CK(clk), .RN(rst_n), .Q(
        y_out_sum0[4]) );
  DFFRHQX1 reg_length6_reg_2_ ( .D(n3620), .CK(clk), .RN(rst_n), .Q(
        reg_length6[2]) );
  DFFRHQX1 y_out_sum8_reg_4_ ( .D(n3556), .CK(clk), .RN(rst_n), .Q(
        y_out_sum8[4]) );
  DFFRHQX1 next_reg_5_ ( .D(n4005), .CK(clk), .RN(rst_n), .Q(next[5]) );
  DFFRHQX1 shift_reg_0_ ( .D(N8752), .CK(clk), .RN(rst_n), .Q(shift[0]) );
  DFFRHQX1 y_out_sum14_reg_4_ ( .D(n3226), .CK(clk), .RN(rst_n), .Q(
        y_out_sum14[4]) );
  DFFRHQX1 shift_reg_1_ ( .D(N8753), .CK(clk), .RN(rst_n), .Q(shift[1]) );
  DFFRHQX1 next_reg_7_ ( .D(n4003), .CK(clk), .RN(rst_n), .Q(next[7]) );
  DFFRHQX1 shift_reg_5_ ( .D(N8757), .CK(clk), .RN(rst_n), .Q(shift[5]) );
  DFFRHQX1 y_out_sum6_reg_4_ ( .D(n3666), .CK(clk), .RN(rst_n), .Q(
        y_out_sum6[4]) );
  DFFRHQX1 reg_length4_reg_2_ ( .D(n3730), .CK(clk), .RN(rst_n), .Q(
        reg_length4[2]) );
  DFFRHQX1 shift_reg_2_ ( .D(N8754), .CK(clk), .RN(rst_n), .Q(shift[2]) );
  DFFRHQX1 reg_length5_reg_1_ ( .D(n3676), .CK(clk), .RN(rst_n), .Q(
        reg_length5[1]) );
  DFFRHQX1 shift_reg_4_ ( .D(N8756), .CK(clk), .RN(rst_n), .Q(shift[4]) );
  DFFRHQX1 y_out_sum2_reg_4_ ( .D(n3886), .CK(clk), .RN(rst_n), .Q(
        y_out_sum2[4]) );
  DFFRHQX1 shift_reg_3_ ( .D(N8755), .CK(clk), .RN(rst_n), .Q(shift[3]) );
  DFFRHQX1 next_reg_6_ ( .D(n4004), .CK(clk), .RN(rst_n), .Q(next[6]) );
  DFFRHQX1 y_out_sum12_reg_4_ ( .D(n3336), .CK(clk), .RN(rst_n), .Q(
        y_out_sum12[4]) );
  DFFRHQX1 y_out_sum10_reg_4_ ( .D(n3446), .CK(clk), .RN(rst_n), .Q(
        y_out_sum10[4]) );
  DFFRHQX1 y_out_sum9_reg_4_ ( .D(n3501), .CK(clk), .RN(rst_n), .Q(
        y_out_sum9[4]) );
  DFFRX1 reg_length14_reg_0_ ( .D(n3182), .CK(clk), .RN(rst_n), .Q(
        reg_length14[0]), .QN(n4952) );
  DFFRHQX1 y_out_sum11_reg_4_ ( .D(n3391), .CK(clk), .RN(rst_n), .Q(
        y_out_sum11[4]) );
  DFFRHQX1 y_out_sum5_reg_3_ ( .D(n3722), .CK(clk), .RN(rst_n), .Q(
        y_out_sum5[3]) );
  DFFRHQX1 y_out_sum1_reg_4_ ( .D(n3932), .CK(clk), .RN(rst_n), .Q(
        y_out_sum1[4]) );
  DFFRHQX1 y_out_sum4_reg_4_ ( .D(n3776), .CK(clk), .RN(rst_n), .Q(
        y_out_sum4[4]) );
  DFFRHQX1 y_out_sum7_reg_4_ ( .D(n3611), .CK(clk), .RN(rst_n), .Q(
        y_out_sum7[4]) );
  DFFRHQX1 y_out_sum0_reg_3_ ( .D(n3973), .CK(clk), .RN(rst_n), .Q(
        y_out_sum0[3]) );
  DFFRHQX1 y_out_sum13_reg_4_ ( .D(n3281), .CK(clk), .RN(rst_n), .Q(
        y_out_sum13[4]) );
  DFFRX1 y_out_sum8_reg_3_ ( .D(n3557), .CK(clk), .RN(rst_n), .Q(y_out_sum8[3]), .QN(n4863) );
  DFFRHQX1 y_out_sum4_reg_3_ ( .D(n3777), .CK(clk), .RN(rst_n), .Q(
        y_out_sum4[3]) );
  DFFRHQX1 reg_length6_reg_0_ ( .D(n3622), .CK(clk), .RN(rst_n), .Q(
        reg_length6[0]) );
  DFFRHQX1 reg_length6_reg_1_ ( .D(n3621), .CK(clk), .RN(rst_n), .Q(
        reg_length6[1]) );
  DFFRHQX1 y_out_sum2_reg_3_ ( .D(n3887), .CK(clk), .RN(rst_n), .Q(
        y_out_sum2[3]) );
  DFFRHQX1 y_out_sum5_reg_2_ ( .D(n3723), .CK(clk), .RN(rst_n), .Q(
        y_out_sum5[2]) );
  DFFRHQX1 reg_length4_reg_0_ ( .D(n3732), .CK(clk), .RN(rst_n), .Q(
        reg_length4[0]) );
  DFFRHQX1 reg_length4_reg_1_ ( .D(n3731), .CK(clk), .RN(rst_n), .Q(
        reg_length4[1]) );
  DFFRHQX1 y_out_sum6_reg_3_ ( .D(n3667), .CK(clk), .RN(rst_n), .Q(
        y_out_sum6[3]) );
  DFFRHQX1 y_out_sum3_reg_3_ ( .D(n3832), .CK(clk), .RN(rst_n), .Q(
        y_out_sum3[3]) );
  DFFRX1 y_out_sum9_reg_3_ ( .D(n3502), .CK(clk), .RN(rst_n), .Q(y_out_sum9[3]), .QN(n4877) );
  DFFRHQX1 y_out_sum1_reg_3_ ( .D(n3933), .CK(clk), .RN(rst_n), .Q(
        y_out_sum1[3]) );
  DFFRX1 reg_length5_reg_0_ ( .D(n3677), .CK(clk), .RN(rst_n), .Q(
        reg_length5[0]), .QN(n4934) );
  DFFRHQX1 current_state_reg_0_ ( .D(next_state[0]), .CK(clk), .RN(rst_n), .Q(
        current_state[0]) );
  DFFRHQX1 current_state_reg_1_ ( .D(next_state[1]), .CK(clk), .RN(rst_n), .Q(
        current_state[1]) );
  DFFRHQX1 y_out_sum4_reg_2_ ( .D(n3778), .CK(clk), .RN(rst_n), .Q(
        y_out_sum4[2]) );
  DFFRX1 y_out_sum14_reg_3_ ( .D(n3227), .CK(clk), .RN(rst_n), .Q(
        y_out_sum14[3]), .QN(n4858) );
  DFFRHQX1 y_out_sum0_reg_2_ ( .D(n3974), .CK(clk), .RN(rst_n), .Q(
        y_out_sum0[2]) );
  DFFRHQX1 y_out_sum6_reg_2_ ( .D(n3668), .CK(clk), .RN(rst_n), .Q(
        y_out_sum6[2]) );
  DFFRHQX1 y_out_sum3_reg_2_ ( .D(n3833), .CK(clk), .RN(rst_n), .Q(
        y_out_sum3[2]) );
  DFFRX1 y_out_sum12_reg_3_ ( .D(n3337), .CK(clk), .RN(rst_n), .Q(
        y_out_sum12[3]), .QN(n4887) );
  DFFRX1 y_out_sum11_reg_3_ ( .D(n3392), .CK(clk), .RN(rst_n), .Q(
        y_out_sum11[3]), .QN(n4853) );
  DFFRX1 y_out_sum8_reg_2_ ( .D(n3558), .CK(clk), .RN(rst_n), .Q(y_out_sum8[2]), .QN(n4913) );
  DFFRHQX1 y_out_sum2_reg_2_ ( .D(n3888), .CK(clk), .RN(rst_n), .Q(
        y_out_sum2[2]) );
  DFFRX1 y_out_sum10_reg_3_ ( .D(n3447), .CK(clk), .RN(rst_n), .Q(
        y_out_sum10[3]), .QN(n4870) );
  DFFRX1 y_out_sum13_reg_3_ ( .D(n3282), .CK(clk), .RN(rst_n), .Q(
        y_out_sum13[3]), .QN(n4880) );
  DFFRHQX1 y_out_sum2_reg_0_ ( .D(n3890), .CK(clk), .RN(rst_n), .Q(
        y_out_sum2[0]) );
  DFFRHQX1 y_out_sum1_reg_2_ ( .D(n3934), .CK(clk), .RN(rst_n), .Q(
        y_out_sum1[2]) );
  DFFRX1 y_out_sum14_reg_2_ ( .D(n3228), .CK(clk), .RN(rst_n), .Q(
        y_out_sum14[2]), .QN(n4906) );
  DFFRX1 y_out_sum10_reg_2_ ( .D(n3448), .CK(clk), .RN(rst_n), .Q(
        y_out_sum10[2]), .QN(n4920) );
  DFFRX1 y_out_sum7_reg_3_ ( .D(n3612), .CK(clk), .RN(rst_n), .Q(y_out_sum7[3]), .QN(n4869) );
  DFFRHQX1 y_out_sum4_reg_0_ ( .D(n3780), .CK(clk), .RN(rst_n), .Q(
        y_out_sum4[0]) );
  DFFRHQX1 y_out_sum14_reg_0_ ( .D(n3230), .CK(clk), .RN(rst_n), .Q(
        y_out_sum14[0]) );
  DFFRX1 y_out_sum9_reg_2_ ( .D(n3503), .CK(clk), .RN(rst_n), .Q(y_out_sum9[2]), .QN(n4922) );
  DFFRX1 y_out_sum12_reg_2_ ( .D(n3338), .CK(clk), .RN(rst_n), .Q(
        y_out_sum12[2]), .QN(n4933) );
  DFFRHQX1 y_out_sum5_reg_0_ ( .D(n3725), .CK(clk), .RN(rst_n), .Q(
        y_out_sum5[0]) );
  DFFRHQX1 y_out_sum9_reg_0_ ( .D(n3505), .CK(clk), .RN(rst_n), .Q(
        y_out_sum9[0]) );
  DFFRHQX1 y_out_sum6_reg_0_ ( .D(n3670), .CK(clk), .RN(rst_n), .Q(
        y_out_sum6[0]) );
  DFFRHQX1 y_out_sum2_reg_1_ ( .D(n3889), .CK(clk), .RN(rst_n), .Q(
        y_out_sum2[1]) );
  DFFRX1 y_out_sum11_reg_2_ ( .D(n3393), .CK(clk), .RN(rst_n), .Q(
        y_out_sum11[2]), .QN(n4903) );
  DFFRHQX1 y_out_sum13_reg_0_ ( .D(n3285), .CK(clk), .RN(rst_n), .Q(
        y_out_sum13[0]) );
  DFFRHQX1 y_out_sum11_reg_0_ ( .D(n3395), .CK(clk), .RN(rst_n), .Q(
        y_out_sum11[0]) );
  DFFRHQX1 y_out_sum12_reg_0_ ( .D(n3340), .CK(clk), .RN(rst_n), .Q(
        y_out_sum12[0]) );
  DFFRHQX1 y_out_sum8_reg_0_ ( .D(n3560), .CK(clk), .RN(rst_n), .Q(
        y_out_sum8[0]) );
  DFFRHQX1 y_out_sum4_reg_1_ ( .D(n3779), .CK(clk), .RN(rst_n), .Q(
        y_out_sum4[1]) );
  DFFRHQX1 y_out_sum10_reg_0_ ( .D(n3450), .CK(clk), .RN(rst_n), .Q(
        y_out_sum10[0]) );
  DFFRHQX1 y_out_sum0_reg_0_ ( .D(n3976), .CK(clk), .RN(rst_n), .Q(
        y_out_sum0[0]) );
  DFFRX1 y_out_sum13_reg_2_ ( .D(n3283), .CK(clk), .RN(rst_n), .Q(
        y_out_sum13[2]), .QN(n4927) );
  DFFRHQX1 y_out_sum14_reg_1_ ( .D(n3229), .CK(clk), .RN(rst_n), .Q(
        y_out_sum14[1]) );
  DFFRHQX1 y_out_sum5_reg_1_ ( .D(n3724), .CK(clk), .RN(rst_n), .Q(
        y_out_sum5[1]) );
  DFFRHQX1 y_out_sum3_reg_0_ ( .D(n3835), .CK(clk), .RN(rst_n), .Q(
        y_out_sum3[0]) );
  DFFRHQX1 y_out_sum6_reg_1_ ( .D(n3669), .CK(clk), .RN(rst_n), .Q(
        y_out_sum6[1]) );
  DFFRHQX1 y_out_sum9_reg_1_ ( .D(n3504), .CK(clk), .RN(rst_n), .Q(
        y_out_sum9[1]) );
  DFFRHQX1 y_out_sum0_reg_1_ ( .D(n3975), .CK(clk), .RN(rst_n), .Q(
        y_out_sum0[1]) );
  DFFRHQX1 y_out_sum11_reg_1_ ( .D(n3394), .CK(clk), .RN(rst_n), .Q(
        y_out_sum11[1]) );
  DFFRHQX1 y_out_sum1_reg_0_ ( .D(n3936), .CK(clk), .RN(rst_n), .Q(
        y_out_sum1[0]) );
  DFFRHQX1 y_out_sum12_reg_1_ ( .D(n3339), .CK(clk), .RN(rst_n), .Q(
        y_out_sum12[1]) );
  DFFRHQX1 y_out_sum8_reg_1_ ( .D(n3559), .CK(clk), .RN(rst_n), .Q(
        y_out_sum8[1]) );
  DFFRHQX1 y_out_sum10_reg_1_ ( .D(n3449), .CK(clk), .RN(rst_n), .Q(
        y_out_sum10[1]) );
  DFFRHQX1 y_out_sum7_reg_0_ ( .D(n3615), .CK(clk), .RN(rst_n), .Q(
        y_out_sum7[0]) );
  DFFRX1 y_out_sum7_reg_2_ ( .D(n3613), .CK(clk), .RN(rst_n), .Q(y_out_sum7[2]), .QN(n4918) );
  DFFRHQX1 y_out_sum3_reg_1_ ( .D(n3834), .CK(clk), .RN(rst_n), .Q(
        y_out_sum3[1]) );
  DFFRHQX1 y_out_sum1_reg_1_ ( .D(n3935), .CK(clk), .RN(rst_n), .Q(
        y_out_sum1[1]) );
  DFFRHQX1 y_out_sum13_reg_1_ ( .D(n3284), .CK(clk), .RN(rst_n), .Q(
        y_out_sum13[1]) );
  DFFRHQX1 y_out_sum7_reg_1_ ( .D(n3614), .CK(clk), .RN(rst_n), .Q(
        y_out_sum7[1]) );
  DFFRHQX1 reg_matrix_size_reg_1_ ( .D(n2850), .CK(clk), .RN(rst_n), .Q(
        reg_matrix_size[1]) );
  DFFSHQX1 reg_matrix_size_reg_3_ ( .D(n2852), .CK(clk), .SN(rst_n), .Q(
        reg_matrix_size[3]) );
  DFFRHQX1 reg_matrix_size_reg_2_ ( .D(n7169), .CK(clk), .RN(rst_n), .Q(
        reg_matrix_size[2]) );
  DFFRHQX1 reg_invalid2_reg_2_ ( .D(n3998), .CK(clk), .RN(rst_n), .Q(
        reg_invalid2[2]) );
  DFFRHQX1 reg_invalid2_reg_5_ ( .D(n3995), .CK(clk), .RN(rst_n), .Q(
        reg_invalid2[5]) );
  DFFRHQX1 reg_invalid2_reg_3_ ( .D(n3997), .CK(clk), .RN(rst_n), .Q(
        reg_invalid2[3]) );
  DFFRHQX1 reg_invalid2_reg_0_ ( .D(n3999), .CK(clk), .RN(rst_n), .Q(
        reg_invalid2[0]) );
  DFFRHQX1 reg_invalid2_reg_4_ ( .D(n3996), .CK(clk), .RN(rst_n), .Q(
        reg_invalid2[4]) );
  DFFRHQX1 reg_invalid2_reg_8_ ( .D(n3992), .CK(clk), .RN(rst_n), .Q(
        reg_invalid2[8]) );
  DFFRHQX1 reg_invalid2_reg_1_ ( .D(n4000), .CK(clk), .RN(rst_n), .Q(
        reg_invalid2[1]) );
  DFFRHQX1 reg_invalid2_reg_7_ ( .D(n3993), .CK(clk), .RN(rst_n), .Q(
        reg_invalid2[7]) );
  DFFRHQX1 reg_invalid2_reg_6_ ( .D(n3994), .CK(clk), .RN(rst_n), .Q(
        reg_invalid2[6]) );
  DFFRHQX1 D1_reg_127_ ( .D(N5385), .CK(clk), .RN(rst_n), .Q(D1[127]) );
  DFFRHQX1 D3_reg_15_ ( .D(N5402), .CK(clk), .RN(rst_n), .Q(D3[15]) );
  DFFRHQX1 A1_reg_5_ ( .D(N4783), .CK(clk), .RN(rst_n), .Q(A1[5]) );
  DFFRHQX1 A1_reg_4_ ( .D(N4782), .CK(clk), .RN(rst_n), .Q(A1[4]) );
  DFFRHQX1 A1_reg_3_ ( .D(N4781), .CK(clk), .RN(rst_n), .Q(A1[3]) );
  DFFRHQX1 A1_reg_2_ ( .D(N4780), .CK(clk), .RN(rst_n), .Q(A1[2]) );
  DFFRHQX1 A1_reg_1_ ( .D(N4779), .CK(clk), .RN(rst_n), .Q(A1[1]) );
  DFFRHQX1 A1_reg_6_ ( .D(N4784), .CK(clk), .RN(rst_n), .Q(A1[6]) );
  DFFRHQX1 A1_reg_0_ ( .D(N4778), .CK(clk), .RN(rst_n), .Q(A1[0]) );
  DFFRXL reg_length00_reg_2_ ( .D(n3174), .CK(clk), .RN(rst_n), .Q(n2841) );
  DFFRXL reg_length00_reg_1_ ( .D(n3175), .CK(clk), .RN(rst_n), .Q(n2840) );
  DFFRHQXL y_out_sum12_reg_25_ ( .D(n3315), .CK(clk), .RN(rst_n), .Q(
        y_out_sum12[25]) );
  DFFRHQXL y_out_sum12_reg_24_ ( .D(n3316), .CK(clk), .RN(rst_n), .Q(
        y_out_sum12[24]) );
  DFFRHQXL y_out_sum7_reg_25_ ( .D(n3590), .CK(clk), .RN(rst_n), .Q(
        y_out_sum7[25]) );
  DFFRHQXL y_out_sum10_reg_25_ ( .D(n3425), .CK(clk), .RN(rst_n), .Q(
        y_out_sum10[25]) );
  DFFRXL y_out_sum12_reg_26_ ( .D(n3314), .CK(clk), .RN(rst_n), .Q(
        y_out_sum12[26]), .QN(n6462) );
  DFFRHQXL y_out_sum7_reg_24_ ( .D(n3591), .CK(clk), .RN(rst_n), .Q(
        y_out_sum7[24]) );
  DFFRHQXL y_out_sum10_reg_24_ ( .D(n3426), .CK(clk), .RN(rst_n), .Q(
        y_out_sum10[24]) );
  DFFRHQXL y_out_sum0_reg_25_ ( .D(n3951), .CK(clk), .RN(rst_n), .Q(
        y_out_sum0[25]) );
  DFFRXL y_out_sum13_reg_26_ ( .D(n3259), .CK(clk), .RN(rst_n), .Q(
        y_out_sum13[26]), .QN(n6408) );
  DFFRXL y_out_sum9_reg_22_ ( .D(n3483), .CK(clk), .RN(rst_n), .Q(
        y_out_sum9[22]), .QN(n6632) );
  DFFRXL y_out_sum9_reg_26_ ( .D(n3479), .CK(clk), .RN(rst_n), .Q(
        y_out_sum9[26]), .QN(n6626) );
  DFFRHQXL y_out_sum0_reg_24_ ( .D(n3952), .CK(clk), .RN(rst_n), .Q(
        y_out_sum0[24]) );
  DFFRXL y_out_sum10_reg_22_ ( .D(n3428), .CK(clk), .RN(rst_n), .Q(
        y_out_sum10[22]), .QN(n6576) );
  DFFRHQXL y_out_sum0_reg_23_ ( .D(n3953), .CK(clk), .RN(rst_n), .Q(
        y_out_sum0[23]) );
  DFFRXL y_out_sum9_reg_23_ ( .D(n3482), .CK(clk), .RN(rst_n), .Q(
        y_out_sum9[23]), .QN(n6630) );
  DFFRXL y_out_sum7_reg_23_ ( .D(n3592), .CK(clk), .RN(rst_n), .Q(
        y_out_sum7[23]), .QN(n6741) );
  DFFRXL y_out_sum10_reg_23_ ( .D(n3427), .CK(clk), .RN(rst_n), .Q(
        y_out_sum10[23]), .QN(n6574) );
  DFFRHQXL y_out_sum0_reg_22_ ( .D(n3954), .CK(clk), .RN(rst_n), .Q(
        y_out_sum0[22]) );
  DFFRHQXL y_out_sum2_reg_25_ ( .D(n3865), .CK(clk), .RN(rst_n), .Q(
        y_out_sum2[25]) );
  DFFRXL y_out_sum8_reg_26_ ( .D(n3534), .CK(clk), .RN(rst_n), .Q(
        y_out_sum8[26]), .QN(n6682) );
  DFFRHQXL y_out_sum14_reg_25_ ( .D(n3205), .CK(clk), .RN(rst_n), .Q(
        y_out_sum14[25]) );
  DFFRHQXL y_out_sum14_reg_24_ ( .D(n3206), .CK(clk), .RN(rst_n), .Q(
        y_out_sum14[24]) );
  DFFRHQXL y_out_sum2_reg_24_ ( .D(n3866), .CK(clk), .RN(rst_n), .Q(
        y_out_sum2[24]) );
  DFFRHQXL y_out_sum3_reg_23_ ( .D(n3812), .CK(clk), .RN(rst_n), .Q(
        y_out_sum3[23]) );
  DFFRHQXL y_out_sum11_reg_25_ ( .D(n3370), .CK(clk), .RN(rst_n), .Q(
        y_out_sum11[25]) );
  DFFRHQXL y_out_sum3_reg_22_ ( .D(n3813), .CK(clk), .RN(rst_n), .Q(
        y_out_sum3[22]) );
  DFFRXL y_out_sum8_reg_23_ ( .D(n3537), .CK(clk), .RN(rst_n), .Q(
        y_out_sum8[23]), .QN(n6686) );
  DFFRHQXL y_out_sum11_reg_24_ ( .D(n3371), .CK(clk), .RN(rst_n), .Q(
        y_out_sum11[24]) );
  DFFRHQXL y_out_sum2_reg_23_ ( .D(n3867), .CK(clk), .RN(rst_n), .Q(
        y_out_sum2[23]) );
  DFFRHQXL y_out_sum2_reg_22_ ( .D(n3868), .CK(clk), .RN(rst_n), .Q(
        y_out_sum2[22]) );
  DFFRXL y_out_sum14_reg_26_ ( .D(n3204), .CK(clk), .RN(rst_n), .Q(
        y_out_sum14[26]), .QN(n6354) );
  DFFRHQXL y_out_sum5_reg_25_ ( .D(n3700), .CK(clk), .RN(rst_n), .Q(
        y_out_sum5[25]) );
  DFFRHQXL y_out_sum1_reg_26_ ( .D(n3910), .CK(clk), .RN(rst_n), .Q(
        y_out_sum1[26]) );
  DFFRXL y_out_sum11_reg_22_ ( .D(n3373), .CK(clk), .RN(rst_n), .Q(
        y_out_sum11[22]), .QN(n6520) );
  DFFRHQXL y_out_sum1_reg_23_ ( .D(n3913), .CK(clk), .RN(rst_n), .Q(
        y_out_sum1[23]) );
  DFFRHQXL y_out_sum1_reg_22_ ( .D(n3914), .CK(clk), .RN(rst_n), .Q(
        y_out_sum1[22]) );
  DFFRHQXL y_out_sum5_reg_24_ ( .D(n3701), .CK(clk), .RN(rst_n), .Q(
        y_out_sum5[24]) );
  DFFRHQXL y_out_sum5_reg_26_ ( .D(n3699), .CK(clk), .RN(rst_n), .Q(
        y_out_sum5[26]) );
  DFFRHQXL y_out_sum5_reg_23_ ( .D(n3702), .CK(clk), .RN(rst_n), .Q(
        y_out_sum5[23]) );
  DFFRXL y_out_sum11_reg_23_ ( .D(n3372), .CK(clk), .RN(rst_n), .Q(
        y_out_sum11[23]), .QN(n6518) );
  DFFRHQXL y_out_sum5_reg_22_ ( .D(n3703), .CK(clk), .RN(rst_n), .Q(
        y_out_sum5[22]) );
  DFFRHQXL y_out_sum6_reg_25_ ( .D(n3645), .CK(clk), .RN(rst_n), .Q(
        y_out_sum6[25]) );
  DFFRHQXL y_out_sum6_reg_24_ ( .D(n3646), .CK(clk), .RN(rst_n), .Q(
        y_out_sum6[24]) );
  DFFRHQXL y_out_sum4_reg_25_ ( .D(n3755), .CK(clk), .RN(rst_n), .Q(
        y_out_sum4[25]) );
  DFFRHQXL y_out_sum4_reg_24_ ( .D(n3756), .CK(clk), .RN(rst_n), .Q(
        y_out_sum4[24]) );
  DFFRHQXL y_out_sum6_reg_23_ ( .D(n3647), .CK(clk), .RN(rst_n), .Q(
        y_out_sum6[23]) );
  DFFRHQXL y_out_sum4_reg_26_ ( .D(n3754), .CK(clk), .RN(rst_n), .Q(
        y_out_sum4[26]) );
  DFFRHQXL y_out_sum6_reg_22_ ( .D(n3648), .CK(clk), .RN(rst_n), .Q(
        y_out_sum6[22]) );
  DFFRHQXL y_out_sum4_reg_23_ ( .D(n3757), .CK(clk), .RN(rst_n), .Q(
        y_out_sum4[23]) );
  DFFRHQXL y_out_sum4_reg_22_ ( .D(n3758), .CK(clk), .RN(rst_n), .Q(
        y_out_sum4[22]) );
  DFFRHQXL reg_length0_reg_1_ ( .D(n3987), .CK(clk), .RN(rst_n), .Q(
        reg_length0[1]) );
  DFFRHQX1 reg_length0_reg_2_ ( .D(n3988), .CK(clk), .RN(rst_n), .Q(
        reg_length0[2]) );
  DFFHQX1 x_in0_reg_0_ ( .D(n2860), .CK(clk), .Q(x_in0[0]) );
  DFFHQX2 x_in7_reg_0_ ( .D(n2986), .CK(clk), .Q(x_in7[0]) );
  DFFHQX2 x_in2_reg_0_ ( .D(n2907), .CK(clk), .Q(x_in2[0]) );
  DFFHQX2 x_in3_reg_0_ ( .D(n2923), .CK(clk), .Q(x_in3[0]) );
  DFFHQX2 x_in6_reg_0_ ( .D(n4029), .CK(clk), .Q(x_in6[0]) );
  DFFHQX2 x_in7_reg_6_ ( .D(n2980), .CK(clk), .Q(x_in7[6]) );
  DFFHQX2 x_in7_reg_5_ ( .D(n2981), .CK(clk), .Q(x_in7[5]) );
  DFFHQX2 x_in7_reg_1_ ( .D(n2985), .CK(clk), .Q(x_in7[1]) );
  DFFHQX2 x_in7_reg_12_ ( .D(n2974), .CK(clk), .Q(x_in7[12]) );
  DFFHQX2 x_in5_reg_8_ ( .D(n2947), .CK(clk), .Q(x_in5[8]) );
  DFFHQX2 x_in5_reg_7_ ( .D(n2948), .CK(clk), .Q(x_in5[7]) );
  DFFHQX2 x_in5_reg_6_ ( .D(n2949), .CK(clk), .Q(x_in5[6]) );
  DFFHQX2 x_in5_reg_5_ ( .D(n2950), .CK(clk), .Q(x_in5[5]) );
  DFFHQX1 x_in5_reg_2_ ( .D(n2953), .CK(clk), .Q(x_in5[2]) );
  DFFHQX2 x_in5_reg_1_ ( .D(n2954), .CK(clk), .Q(x_in5[1]) );
  DFFHQX2 x_in5_reg_14_ ( .D(n2941), .CK(clk), .Q(x_in5[14]) );
  DFFHQX2 x_in5_reg_0_ ( .D(n2955), .CK(clk), .Q(x_in5[0]) );
  DFFHQX2 x_in6_reg_9_ ( .D(n2962), .CK(clk), .Q(x_in6[9]) );
  DFFHQX2 x_in6_reg_5_ ( .D(n2966), .CK(clk), .Q(x_in6[5]) );
  DFFHQX2 x_in6_reg_4_ ( .D(n2967), .CK(clk), .Q(x_in6[4]) );
  DFFHQX2 x_in6_reg_3_ ( .D(n2968), .CK(clk), .Q(x_in6[3]) );
  DFFHQX2 x_in6_reg_12_ ( .D(n2959), .CK(clk), .Q(x_in6[12]) );
  DFFHQX2 x_in6_reg_11_ ( .D(n2960), .CK(clk), .Q(x_in6[11]) );
  DFFHQX2 x_in6_reg_10_ ( .D(n2961), .CK(clk), .Q(x_in6[10]) );
  DFFHQX2 x_in4_reg_5_ ( .D(n2934), .CK(clk), .Q(x_in4[5]) );
  DFFHQX2 x_in4_reg_4_ ( .D(n2935), .CK(clk), .Q(x_in4[4]) );
  DFFHQX2 x_in4_reg_3_ ( .D(n2936), .CK(clk), .Q(x_in4[3]) );
  DFFHQX2 x_in4_reg_1_ ( .D(n2938), .CK(clk), .Q(x_in4[1]) );
  DFFHQX2 x_in4_reg_10_ ( .D(n2929), .CK(clk), .Q(x_in4[10]) );
  DFFHQX2 x_in4_reg_0_ ( .D(n2939), .CK(clk), .Q(x_in4[0]) );
  DFFHQX2 x_in3_reg_9_ ( .D(n2914), .CK(clk), .Q(x_in3[9]) );
  DFFHQX2 x_in3_reg_8_ ( .D(n2915), .CK(clk), .Q(x_in3[8]) );
  DFFHQX2 x_in3_reg_6_ ( .D(n2917), .CK(clk), .Q(x_in3[6]) );
  DFFHQX1 x_in3_reg_5_ ( .D(n2918), .CK(clk), .Q(x_in3[5]) );
  DFFHQX1 x_in3_reg_4_ ( .D(n2919), .CK(clk), .Q(x_in3[4]) );
  DFFHQX1 x_in3_reg_3_ ( .D(n2920), .CK(clk), .Q(x_in3[3]) );
  DFFHQX2 x_in3_reg_1_ ( .D(n2922), .CK(clk), .Q(x_in3[1]) );
  DFFHQX1 x_in3_reg_14_ ( .D(n2909), .CK(clk), .Q(x_in3[14]) );
  DFFHQX2 x_in3_reg_10_ ( .D(n2913), .CK(clk), .Q(x_in3[10]) );
  DFFHQX2 x_in2_reg_9_ ( .D(n2898), .CK(clk), .Q(x_in2[9]) );
  DFFHQX1 x_in2_reg_8_ ( .D(n2899), .CK(clk), .Q(x_in2[8]) );
  DFFHQX1 x_in2_reg_7_ ( .D(n2900), .CK(clk), .Q(x_in2[7]) );
  DFFHQX2 x_in2_reg_6_ ( .D(n2901), .CK(clk), .Q(x_in2[6]) );
  DFFHQX2 x_in2_reg_5_ ( .D(n2902), .CK(clk), .Q(x_in2[5]) );
  DFFHQX2 x_in2_reg_4_ ( .D(n2903), .CK(clk), .Q(x_in2[4]) );
  DFFHQX1 x_in2_reg_3_ ( .D(n2904), .CK(clk), .Q(x_in2[3]) );
  DFFHQX1 x_in2_reg_2_ ( .D(n2905), .CK(clk), .Q(x_in2[2]) );
  DFFHQX1 x_in2_reg_1_ ( .D(n2906), .CK(clk), .Q(x_in2[1]) );
  DFFHQX1 x_in2_reg_15_ ( .D(n2892), .CK(clk), .Q(x_in2[15]) );
  DFFHQX1 x_in2_reg_14_ ( .D(n2893), .CK(clk), .Q(x_in2[14]) );
  DFFHQX1 x_in2_reg_13_ ( .D(n2894), .CK(clk), .Q(x_in2[13]) );
  DFFHQX2 x_in2_reg_10_ ( .D(n2897), .CK(clk), .Q(x_in2[10]) );
  DFFHQX2 x_in0_reg_9_ ( .D(n2875), .CK(clk), .Q(x_in0[9]) );
  DFFHQX2 x_in0_reg_8_ ( .D(n2874), .CK(clk), .Q(x_in0[8]) );
  DFFHQX2 x_in0_reg_7_ ( .D(n2873), .CK(clk), .Q(x_in0[7]) );
  DFFHQX2 x_in0_reg_6_ ( .D(n2872), .CK(clk), .Q(x_in0[6]) );
  DFFHQX2 x_in0_reg_5_ ( .D(n2871), .CK(clk), .Q(x_in0[5]) );
  DFFHQX1 x_in0_reg_4_ ( .D(n2870), .CK(clk), .Q(x_in0[4]) );
  DFFHQX1 x_in0_reg_3_ ( .D(n2869), .CK(clk), .Q(x_in0[3]) );
  DFFHQX1 x_in0_reg_2_ ( .D(n2868), .CK(clk), .Q(x_in0[2]) );
  DFFHQX1 x_in0_reg_1_ ( .D(n2867), .CK(clk), .Q(x_in0[1]) );
  DFFHQX1 x_in0_reg_15_ ( .D(n2866), .CK(clk), .Q(x_in0[15]) );
  DFFHQX1 x_in0_reg_14_ ( .D(n2865), .CK(clk), .Q(x_in0[14]) );
  DFFHQX1 x_in0_reg_13_ ( .D(n2864), .CK(clk), .Q(x_in0[13]) );
  DFFHQX2 x_in0_reg_12_ ( .D(n2863), .CK(clk), .Q(x_in0[12]) );
  DFFHQX2 x_in0_reg_11_ ( .D(n2862), .CK(clk), .Q(x_in0[11]) );
  DFFHQX2 x_in0_reg_10_ ( .D(n2861), .CK(clk), .Q(x_in0[10]) );
  DFFHQX2 x_in1_reg_9_ ( .D(n2891), .CK(clk), .Q(x_in1[9]) );
  DFFHQX2 x_in1_reg_8_ ( .D(n2890), .CK(clk), .Q(x_in1[8]) );
  DFFHQX2 x_in1_reg_7_ ( .D(n2889), .CK(clk), .Q(x_in1[7]) );
  DFFHQX1 x_in1_reg_4_ ( .D(n2886), .CK(clk), .Q(x_in1[4]) );
  DFFHQX1 x_in1_reg_3_ ( .D(n2885), .CK(clk), .Q(x_in1[3]) );
  DFFHQX2 x_in1_reg_2_ ( .D(n2884), .CK(clk), .Q(x_in1[2]) );
  DFFHQX1 x_in1_reg_1_ ( .D(n2883), .CK(clk), .Q(x_in1[1]) );
  DFFHQX1 x_in1_reg_15_ ( .D(n2882), .CK(clk), .Q(x_in1[15]) );
  DFFHQX2 x_in1_reg_14_ ( .D(n2881), .CK(clk), .Q(x_in1[14]) );
  DFFHQX1 x_in1_reg_13_ ( .D(n2880), .CK(clk), .Q(x_in1[13]) );
  DFFHQX1 x_in1_reg_12_ ( .D(n2879), .CK(clk), .Q(x_in1[12]) );
  DFFHQX2 x_in1_reg_10_ ( .D(n2877), .CK(clk), .Q(x_in1[10]) );
  DFFHQX2 x_in1_reg_0_ ( .D(n2876), .CK(clk), .Q(x_in1[0]) );
  DFFHQX2 w_in7_reg_8_ ( .D(n7137), .CK(clk), .Q(w_in7[8]) );
  DFFHQX2 w_in3_reg_8_ ( .D(n3010), .CK(clk), .Q(w_in3[8]) );
  DFFHQX2 w_in7_reg_6_ ( .D(n7139), .CK(clk), .Q(w_in7[6]) );
  DFFHQX2 w_in3_reg_6_ ( .D(n3012), .CK(clk), .Q(w_in3[6]) );
  DFFHQX1 w_in4_reg_15_ ( .D(n3099), .CK(clk), .Q(w_in4[15]) );
  DFFHQX1 w_in4_reg_14_ ( .D(n3100), .CK(clk), .Q(w_in4[14]) );
  DFFHQX1 w_in4_reg_13_ ( .D(n3101), .CK(clk), .Q(w_in4[13]) );
  DFFHQX2 w_in4_reg_12_ ( .D(n3102), .CK(clk), .Q(w_in4[12]) );
  DFFHQX2 w_in4_reg_11_ ( .D(n3103), .CK(clk), .Q(w_in4[11]) );
  DFFHQX2 w_in4_reg_10_ ( .D(n3104), .CK(clk), .Q(w_in4[10]) );
  DFFHQX2 w_in4_reg_9_ ( .D(n3105), .CK(clk), .Q(w_in4[9]) );
  DFFHQX2 w_in4_reg_8_ ( .D(n3106), .CK(clk), .Q(w_in4[8]) );
  DFFHQX2 w_in4_reg_6_ ( .D(n3108), .CK(clk), .Q(w_in4[6]) );
  DFFHQX2 w_in4_reg_4_ ( .D(n3110), .CK(clk), .Q(w_in4[4]) );
  DFFHQX2 w_in4_reg_2_ ( .D(n3112), .CK(clk), .Q(w_in4[2]) );
  DFFHQX2 w_in7_reg_4_ ( .D(n7141), .CK(clk), .Q(w_in7[4]) );
  DFFHQX2 w_in3_reg_4_ ( .D(n3014), .CK(clk), .Q(w_in3[4]) );
  DFFHQX2 w_in4_reg_0_ ( .D(n3114), .CK(clk), .Q(w_in4[0]) );
  DFFHQX1 w_in5_reg_15_ ( .D(n3083), .CK(clk), .Q(w_in5[15]) );
  DFFHQX2 w_in5_reg_13_ ( .D(n3085), .CK(clk), .Q(w_in5[13]) );
  DFFHQX2 w_in5_reg_12_ ( .D(n3086), .CK(clk), .Q(w_in5[12]) );
  DFFHQX2 w_in5_reg_11_ ( .D(n3087), .CK(clk), .Q(w_in5[11]) );
  DFFHQX2 w_in5_reg_10_ ( .D(n3088), .CK(clk), .Q(w_in5[10]) );
  DFFHQX2 w_in5_reg_9_ ( .D(n3089), .CK(clk), .Q(w_in5[9]) );
  DFFHQX2 w_in5_reg_8_ ( .D(n3090), .CK(clk), .Q(w_in5[8]) );
  DFFHQX2 w_in5_reg_7_ ( .D(n3091), .CK(clk), .Q(w_in5[7]) );
  DFFHQX2 w_in5_reg_6_ ( .D(n3092), .CK(clk), .Q(w_in5[6]) );
  DFFHQX2 w_in1_reg_3_ ( .D(n3031), .CK(clk), .Q(w_in1[3]) );
  DFFHQX1 w_in5_reg_0_ ( .D(n3098), .CK(clk), .Q(w_in5[0]) );
  DFFHQX1 w_in6_reg_15_ ( .D(n7143), .CK(clk), .Q(w_in6[15]) );
  DFFHQX1 w_in2_reg_15_ ( .D(n3067), .CK(clk), .Q(w_in2[15]) );
  DFFHQX2 w_in7_reg_2_ ( .D(n7145), .CK(clk), .Q(w_in7[2]) );
  DFFHQX2 w_in1_reg_2_ ( .D(n3032), .CK(clk), .Q(w_in1[2]) );
  DFFHQX2 w_in3_reg_2_ ( .D(n3016), .CK(clk), .Q(w_in3[2]) );
  DFFHQX2 w_in6_reg_13_ ( .D(n7146), .CK(clk), .Q(w_in6[13]) );
  DFFHQX2 w_in6_reg_12_ ( .D(n7147), .CK(clk), .Q(w_in6[12]) );
  DFFHQX2 w_in2_reg_12_ ( .D(n3070), .CK(clk), .Q(w_in2[12]) );
  DFFHQX1 w_in6_reg_10_ ( .D(n7149), .CK(clk), .Q(w_in6[10]) );
  DFFHQX2 w_in2_reg_10_ ( .D(n3072), .CK(clk), .Q(w_in2[10]) );
  DFFHQX2 w_in6_reg_8_ ( .D(n7151), .CK(clk), .Q(w_in6[8]) );
  DFFHQX2 w_in2_reg_8_ ( .D(n3074), .CK(clk), .Q(w_in2[8]) );
  DFFHQX2 w_in6_reg_6_ ( .D(n7153), .CK(clk), .Q(w_in6[6]) );
  DFFHQX2 w_in2_reg_6_ ( .D(n3076), .CK(clk), .Q(w_in2[6]) );
  DFFHQX2 w_in6_reg_4_ ( .D(n7155), .CK(clk), .Q(w_in6[4]) );
  DFFHQX2 w_in2_reg_4_ ( .D(n3078), .CK(clk), .Q(w_in2[4]) );
  DFFHQX2 w_in6_reg_2_ ( .D(n7158), .CK(clk), .Q(w_in6[2]) );
  DFFHQX2 w_in2_reg_2_ ( .D(n3080), .CK(clk), .Q(w_in2[2]) );
  DFFHQX1 w_in6_reg_0_ ( .D(n7160), .CK(clk), .Q(w_in6[0]) );
  DFFHQX2 w_in2_reg_0_ ( .D(n3082), .CK(clk), .Q(w_in2[0]) );
  DFFHQX2 w_in7_reg_15_ ( .D(n7161), .CK(clk), .Q(w_in7[15]) );
  DFFHQX1 w_in3_reg_15_ ( .D(n3003), .CK(clk), .Q(w_in3[15]) );
  DFFHQX2 w_in7_reg_14_ ( .D(n7162), .CK(clk), .Q(w_in7[14]) );
  DFFHQX2 w_in7_reg_13_ ( .D(n7163), .CK(clk), .Q(w_in7[13]) );
  DFFHQX2 w_in7_reg_12_ ( .D(n7164), .CK(clk), .Q(w_in7[12]) );
  DFFHQX1 w_in0_reg_15_ ( .D(n3035), .CK(clk), .Q(w_in0[15]) );
  DFFHQX2 w_in0_reg_14_ ( .D(n3036), .CK(clk), .Q(w_in0[14]) );
  DFFHQX2 w_in0_reg_12_ ( .D(n3038), .CK(clk), .Q(w_in0[12]) );
  DFFHQX2 w_in0_reg_10_ ( .D(n3040), .CK(clk), .Q(w_in0[10]) );
  DFFHQX2 w_in0_reg_8_ ( .D(n3042), .CK(clk), .Q(w_in0[8]) );
  DFFHQX2 w_in7_reg_11_ ( .D(n7165), .CK(clk), .Q(w_in7[11]) );
  DFFHQX2 w_in0_reg_6_ ( .D(n3044), .CK(clk), .Q(w_in0[6]) );
  DFFHQX2 w_in0_reg_4_ ( .D(n3046), .CK(clk), .Q(w_in0[4]) );
  DFFHQX2 w_in0_reg_2_ ( .D(n3048), .CK(clk), .Q(w_in0[2]) );
  DFFHQX1 w_in0_reg_0_ ( .D(n3050), .CK(clk), .Q(w_in0[0]) );
  DFFHQX1 w_in1_reg_15_ ( .D(n3019), .CK(clk), .Q(w_in1[15]) );
  DFFHQX2 w_in1_reg_14_ ( .D(n3020), .CK(clk), .Q(w_in1[14]) );
  DFFHQX2 w_in7_reg_10_ ( .D(n7166), .CK(clk), .Q(w_in7[10]) );
  DFFHQX2 w_in3_reg_10_ ( .D(n3008), .CK(clk), .Q(w_in3[10]) );
  DFFHQX2 w_in1_reg_12_ ( .D(n3022), .CK(clk), .Q(w_in1[12]) );
  DFFHQX1 w_in1_reg_8_ ( .D(n3026), .CK(clk), .Q(w_in1[8]) );
  DFFHQX2 w_in1_reg_5_ ( .D(n3029), .CK(clk), .Q(w_in1[5]) );
  DFFHQX2 w_in7_reg_0_ ( .D(n7167), .CK(clk), .Q(w_in7[0]) );
  DFFHQX2 w_in3_reg_0_ ( .D(n3018), .CK(clk), .Q(w_in3[0]) );
  DFFHQX1 w_in5_reg_2_ ( .D(n3096), .CK(clk), .Q(w_in5[2]) );
  DFFHQX1 w_in5_reg_4_ ( .D(n3094), .CK(clk), .Q(w_in5[4]) );
  DFFTRX2 w_in6_reg_7_ ( .D(1'b1), .RN(n7152), .CK(clk), .Q(w_in6[7]), .QN(
        n5598) );
  DFFHQX4 x_in7_reg_11_ ( .D(n2975), .CK(clk), .Q(x_in7[11]) );
  DFFHQX4 x_in4_reg_14_ ( .D(n2925), .CK(clk), .Q(x_in4[14]) );
  DFFHQX4 x_in6_reg_6_ ( .D(n2965), .CK(clk), .Q(x_in6[6]) );
  DFFHQX4 x_in7_reg_4_ ( .D(n2982), .CK(clk), .Q(x_in7[4]) );
  DFFHQX4 x_in4_reg_13_ ( .D(n2926), .CK(clk), .Q(x_in4[13]) );
  DFFHQX4 x_in7_reg_13_ ( .D(n2973), .CK(clk), .Q(x_in7[13]) );
  DFFHQX4 x_in4_reg_15_ ( .D(n2924), .CK(clk), .Q(x_in4[15]) );
  DFFHQX4 x_in7_reg_10_ ( .D(n2976), .CK(clk), .Q(x_in7[10]) );
  DFFHQX4 x_in4_reg_9_ ( .D(n2930), .CK(clk), .Q(x_in4[9]) );
  DFFHQX4 x_in7_reg_9_ ( .D(n2977), .CK(clk), .Q(x_in7[9]) );
  DFFHQX4 x_in4_reg_12_ ( .D(n2927), .CK(clk), .Q(x_in4[12]) );
  DFFHQX4 x_in4_reg_8_ ( .D(n2931), .CK(clk), .Q(x_in4[8]) );
  DFFHQX4 x_in7_reg_7_ ( .D(n2979), .CK(clk), .Q(x_in7[7]) );
  DFFHQX4 w_in1_reg_10_ ( .D(n3024), .CK(clk), .Q(w_in1[10]) );
  DFFHQX4 x_in7_reg_8_ ( .D(n2978), .CK(clk), .Q(x_in7[8]) );
  DFFHQX4 x_in1_reg_11_ ( .D(n2878), .CK(clk), .Q(x_in1[11]) );
  DFFHQX2 w_in1_reg_4_ ( .D(n3030), .CK(clk), .Q(w_in1[4]) );
  DFFHQX4 x_in4_reg_11_ ( .D(n2928), .CK(clk), .Q(x_in4[11]) );
  DFFHQX4 x_in5_reg_11_ ( .D(n2944), .CK(clk), .Q(x_in5[11]) );
  DFFHQX2 w_in1_reg_6_ ( .D(n3028), .CK(clk), .Q(w_in1[6]) );
  DFFHQX4 x_in5_reg_12_ ( .D(n2943), .CK(clk), .Q(x_in5[12]) );
  DFFHQX4 x_in6_reg_15_ ( .D(n2956), .CK(clk), .Q(x_in6[15]) );
  DFFHQX4 x_in7_reg_3_ ( .D(n2983), .CK(clk), .Q(x_in7[3]) );
  DFFHQX4 x_in7_reg_15_ ( .D(n2971), .CK(clk), .Q(x_in7[15]) );
  DFFHQX4 x_in7_reg_14_ ( .D(n2972), .CK(clk), .Q(x_in7[14]) );
  DFFHQX4 x_in6_reg_1_ ( .D(n2970), .CK(clk), .Q(x_in6[1]) );
  DFFHQX4 x_in5_reg_15_ ( .D(n2940), .CK(clk), .Q(x_in5[15]) );
  DFFHQX2 x_in5_reg_10_ ( .D(n2945), .CK(clk), .Q(x_in5[10]) );
  DFFHQX4 x_in6_reg_14_ ( .D(n2957), .CK(clk), .Q(x_in6[14]) );
  DFFHQX4 x_in5_reg_9_ ( .D(n2946), .CK(clk), .Q(x_in5[9]) );
  DFFHQX2 w_in5_reg_14_ ( .D(n3084), .CK(clk), .Q(w_in5[14]) );
  DFFHQX2 x_in4_reg_2_ ( .D(n2937), .CK(clk), .Q(x_in4[2]) );
  DFFHQX4 x_in1_reg_6_ ( .D(n2888), .CK(clk), .Q(x_in1[6]) );
  DFFHQX4 x_in4_reg_7_ ( .D(n2932), .CK(clk), .Q(x_in4[7]) );
  DFFHQX4 x_in3_reg_12_ ( .D(n2911), .CK(clk), .Q(x_in3[12]) );
  DFFHQX4 x_in6_reg_8_ ( .D(n2963), .CK(clk), .Q(x_in6[8]) );
  DFFHQX4 x_in5_reg_13_ ( .D(n2942), .CK(clk), .Q(x_in5[13]) );
  DFFHQX4 x_in6_reg_13_ ( .D(n2958), .CK(clk), .Q(x_in6[13]) );
  DFFHQX4 x_in3_reg_11_ ( .D(n2912), .CK(clk), .Q(x_in3[11]) );
  DFFHQX2 w_in6_reg_14_ ( .D(n7144), .CK(clk), .Q(w_in6[14]) );
  DFFHQX4 x_in1_reg_5_ ( .D(n2887), .CK(clk), .Q(x_in1[5]) );
  DFFHQX2 x_in6_reg_7_ ( .D(n2964), .CK(clk), .Q(x_in6[7]) );
  DFFHQX2 x_in5_reg_3_ ( .D(n2952), .CK(clk), .Q(x_in5[3]) );
  DFFHQX4 x_in3_reg_7_ ( .D(n2916), .CK(clk), .Q(x_in3[7]) );
  DFFHQX4 x_in2_reg_12_ ( .D(n2895), .CK(clk), .Q(x_in2[12]) );
  DFFHQX4 x_in7_reg_2_ ( .D(n2984), .CK(clk), .Q(x_in7[2]) );
  DFFHQX2 x_in5_reg_4_ ( .D(n2951), .CK(clk), .Q(x_in5[4]) );
  DFFHQX4 x_in3_reg_15_ ( .D(n2908), .CK(clk), .Q(x_in3[15]) );
  DFFHQX4 x_in4_reg_6_ ( .D(n2933), .CK(clk), .Q(x_in4[6]) );
  DFFHQX4 w_in3_reg_12_ ( .D(n3006), .CK(clk), .Q(w_in3[12]) );
  DFFHQX4 w_in3_reg_14_ ( .D(n3004), .CK(clk), .Q(w_in3[14]) );
  DFFHQX4 w_in1_reg_0_ ( .D(n3034), .CK(clk), .Q(w_in1[0]) );
  DFFHQX2 x_in3_reg_13_ ( .D(n2910), .CK(clk), .Q(x_in3[13]) );
  DFFRHQXL y_out_sum3_reg_39_ ( .D(n3836), .CK(clk), .RN(rst_n), .Q(
        y_out_sum3[39]) );
  DFFHQX2 x_in2_reg_11_ ( .D(n2896), .CK(clk), .Q(x_in2[11]) );
  DFFHQX2 x_in3_reg_2_ ( .D(n2921), .CK(clk), .Q(x_in3[2]) );
  DFFHQX2 x_in6_reg_2_ ( .D(n2969), .CK(clk), .Q(x_in6[2]) );
  DFFHQX4 w_in2_reg_14_ ( .D(n3068), .CK(clk), .Q(w_in2[14]) );
  INVX4 U4941 ( .A(n5563), .Y(n5562) );
  INVX4 U4942 ( .A(n5561), .Y(n5559) );
  INVX4 U4943 ( .A(n5494), .Y(n5492) );
  OR2X4 U4944 ( .A(n6006), .B(n6019), .Y(n6026) );
  OR2X4 U4945 ( .A(n5999), .B(n5995), .Y(n6019) );
  INVX4 U4946 ( .A(n5550), .Y(n5549) );
  CLKINVX4 U4947 ( .A(sum[32]), .Y(n5550) );
  CLKINVX3 U4948 ( .A(n5519), .Y(n4986) );
  CLKINVX4 U4949 ( .A(n5519), .Y(n5518) );
  OAI2BB1X2 U4950 ( .A0N(N5845), .A1N(n4990), .B0(n6045), .Y(n3671) );
  CLKINVX4 U4951 ( .A(sum[31]), .Y(n5548) );
  CLKINVX8 U4952 ( .A(n4839), .Y(n4841) );
  OR2X4 U4953 ( .A(n6004), .B(n6000), .Y(n6006) );
  CLKINVX4 U4954 ( .A(sum[37]), .Y(n5561) );
  BUFX8 U4955 ( .A(n5533), .Y(n4846) );
  CLKINVX8 U4956 ( .A(n5550), .Y(n5347) );
  CLKINVX4 U4957 ( .A(n5564), .Y(n4839) );
  INVX2 U4958 ( .A(n4839), .Y(n4840) );
  INVX8 U4959 ( .A(n5548), .Y(n5547) );
  CLKINVX8 U4960 ( .A(n5546), .Y(n5545) );
  INVX3 U4961 ( .A(sum[30]), .Y(n5546) );
  INVX2 U4962 ( .A(sum[1]), .Y(n5478) );
  INVX2 U4963 ( .A(sum[3]), .Y(n5483) );
  INVX2 U4964 ( .A(sum[4]), .Y(n5486) );
  INVX2 U4965 ( .A(sum[29]), .Y(n5544) );
  OR2X1 U4966 ( .A(sum[36]), .B(sum[33]), .Y(n5999) );
  NAND2X1 U4967 ( .A(reg_length0[1]), .B(n7020), .Y(n4981) );
  INVX2 U4968 ( .A(n5528), .Y(n5527) );
  INVX4 U4969 ( .A(n5537), .Y(n5535) );
  BUFX4 U4970 ( .A(n5562), .Y(n4842) );
  INVX2 U4971 ( .A(n5566), .Y(n5564) );
  BUFX8 U4972 ( .A(n5562), .Y(n4843) );
  INVX2 U4973 ( .A(sum[36]), .Y(n5563) );
  NAND2X1 U4974 ( .A(reg_length0[2]), .B(n7022), .Y(n4979) );
  OAI2BB1X1 U4975 ( .A0N(n5955), .A1N(n5558), .B0(n6030), .Y(n6784) );
  INVX2 U4976 ( .A(n5557), .Y(n5555) );
  CLKINVX1 U4977 ( .A(sum[38]), .Y(n5557) );
  BUFX2 U4978 ( .A(n4970), .Y(n4844) );
  CLKINVXL U4979 ( .A(n5512), .Y(n4970) );
  BUFX2 U4980 ( .A(n5533), .Y(n4845) );
  OR2X1 U4981 ( .A(n2788), .B(n6391), .Y(n4847) );
  OR2X1 U4982 ( .A(n102), .B(n2376), .Y(n4848) );
  INVX2 U4983 ( .A(x_in6[0]), .Y(n5469) );
  INVX2 U4984 ( .A(x_in3[0]), .Y(n5472) );
  INVX2 U4985 ( .A(x_in2[0]), .Y(n5473) );
  OR2X1 U4986 ( .A(n2106), .B(n6444), .Y(n4850) );
  OR3X2 U4987 ( .A(n7230), .B(n6552), .C(n2723), .Y(n4851) );
  INVX2 U4988 ( .A(x_in5[0]), .Y(n5470) );
  INVX2 U4989 ( .A(x_in4[0]), .Y(n5471) );
  CLKINVX4 U4990 ( .A(n5512), .Y(n5511) );
  INVX1 U4991 ( .A(sum[22]), .Y(n5528) );
  INVX2 U4992 ( .A(sum[11]), .Y(n5503) );
  INVX4 U4993 ( .A(n5503), .Y(n5502) );
  INVX2 U4994 ( .A(sum[33]), .Y(n5552) );
  INVX2 U4995 ( .A(n5522), .Y(n4983) );
  CLKINVX2 U4996 ( .A(n5522), .Y(n5521) );
  INVX2 U4997 ( .A(sum[18]), .Y(n5519) );
  INVX4 U4998 ( .A(sum[27]), .Y(n5540) );
  INVX4 U4999 ( .A(n5540), .Y(n5538) );
  INVX2 U5000 ( .A(sum[25]), .Y(n5534) );
  INVX2 U5001 ( .A(n5534), .Y(n5533) );
  INVX2 U5002 ( .A(sum[24]), .Y(n5532) );
  INVX4 U5003 ( .A(n5532), .Y(n5531) );
  INVX4 U5004 ( .A(n5496), .Y(n5495) );
  INVX4 U5005 ( .A(n5524), .Y(n5523) );
  INVX2 U5006 ( .A(sum[17]), .Y(n5517) );
  INVX2 U5007 ( .A(sum[9]), .Y(n5498) );
  INVX2 U5008 ( .A(n5542), .Y(n4972) );
  INVX2 U5009 ( .A(n5554), .Y(n5553) );
  INVX2 U5010 ( .A(next[0]), .Y(n5898) );
  INVX2 U5012 ( .A(n5561), .Y(n5560) );
  INVX4 U5013 ( .A(n5498), .Y(n5497) );
  OR2X4 U5014 ( .A(sum[39]), .B(n6026), .Y(n6989) );
  INVX2 U5015 ( .A(sum[15]), .Y(n5512) );
  CLKINVX4 U5016 ( .A(n5510), .Y(n5509) );
  INVX2 U5017 ( .A(sum[14]), .Y(n5510) );
  CLKINVX2 U5018 ( .A(n5488), .Y(n4967) );
  INVX2 U5019 ( .A(sum[5]), .Y(n5488) );
  INVX2 U5020 ( .A(sum[8]), .Y(n5496) );
  INVX2 U5021 ( .A(n5508), .Y(n4968) );
  CLKINVX2 U5022 ( .A(n5508), .Y(n4969) );
  INVX2 U5023 ( .A(sum[13]), .Y(n5508) );
  CLKINVX2 U5024 ( .A(n5491), .Y(n4971) );
  CLKINVX2 U5025 ( .A(n5491), .Y(n5489) );
  INVX2 U5026 ( .A(sum[6]), .Y(n5491) );
  OAI221X2 U5027 ( .A0(n7001), .A1(n7002), .B0(n5350), .B1(n7000), .C0(n6999), 
        .Y(n7010) );
  CLKINVXL U5028 ( .A(n5546), .Y(n4973) );
  CLKINVXL U5029 ( .A(n5546), .Y(n4974) );
  CLKINVX2 U5030 ( .A(n5540), .Y(n4975) );
  CLKINVX2 U5031 ( .A(n5530), .Y(n4976) );
  CLKINVX2 U5032 ( .A(n5530), .Y(n4977) );
  CLKINVX3 U5033 ( .A(n5530), .Y(n5529) );
  INVX4 U5034 ( .A(sum[23]), .Y(n5530) );
  INVX4 U5035 ( .A(n5515), .Y(n5513) );
  CLKINVX3 U5036 ( .A(n5519), .Y(n4985) );
  CLKINVX8 U5037 ( .A(n5552), .Y(n5551) );
  NOR2X1 U5038 ( .A(n2804), .B(n6777), .Y(n5006) );
  CLKINVX2 U5039 ( .A(n5517), .Y(n4978) );
  NAND2X4 U5040 ( .A(n5006), .B(n6989), .Y(n4980) );
  AND3X4 U5041 ( .A(n4979), .B(n4980), .C(n4981), .Y(n6991) );
  AND2X4 U5042 ( .A(n6991), .B(n6990), .Y(n7000) );
  INVX4 U5043 ( .A(n5566), .Y(n5565) );
  CLKINVXL U5044 ( .A(n5546), .Y(n4982) );
  CLKINVX2 U5045 ( .A(n5522), .Y(n5520) );
  CLKINVXL U5046 ( .A(n5566), .Y(n4984) );
  CLKINVX4 U5047 ( .A(sum[35]), .Y(n5566) );
  INVX2 U5048 ( .A(n5483), .Y(n5481) );
  AOI2BB1XL U5049 ( .A0N(n5485), .A1N(n2353), .B0(sum[5]), .Y(n2352) );
  OAI2BB1XL U5050 ( .A0N(N5758), .A1N(n4989), .B0(n6146), .Y(n3746) );
  OAI2BB1XL U5051 ( .A0N(N6497), .A1N(n4993), .B0(n6389), .Y(n3231) );
  OAI2BB1XL U5052 ( .A0N(N5844), .A1N(n4990), .B0(n6046), .Y(n3632) );
  OAI2BB1XL U5053 ( .A0N(N6456), .A1N(n4992), .B0(n6443), .Y(n3286) );
  OAI2BB1XL U5054 ( .A0N(N5762), .A1N(n4989), .B0(n6142), .Y(n3742) );
  OAI2BB1XL U5055 ( .A0N(N5795), .A1N(n4991), .B0(n6102), .Y(n3695) );
  OAI2BB1XL U5056 ( .A0N(N5711), .A1N(n4998), .B0(n6201), .Y(n3807) );
  CLKINVXL U5057 ( .A(n6027), .Y(n5952) );
  OR2X1 U5058 ( .A(n5514), .B(n4844), .Y(n5981) );
  OR2X1 U5059 ( .A(n5505), .B(sum[11]), .Y(n5978) );
  CLKINVXL U5060 ( .A(n5483), .Y(n5482) );
  AOI2BB1X1 U5061 ( .A0N(n2352), .A1N(n5489), .B0(n5493), .Y(n2351) );
  CLKINVXL U5062 ( .A(n6989), .Y(n6036) );
  CLKINVX1 U5063 ( .A(n6011), .Y(n6012) );
  OR2X2 U5064 ( .A(n5556), .B(n5560), .Y(n6004) );
  OR2X2 U5065 ( .A(sum[36]), .B(n5565), .Y(n6000) );
  CLKINVXL U5066 ( .A(n6019), .Y(n6020) );
  OR2XL U5067 ( .A(n4986), .B(n5516), .Y(n5985) );
  OR2XL U5068 ( .A(n5992), .B(n5998), .Y(n6007) );
  OR2XL U5069 ( .A(n5500), .B(sum[9]), .Y(n5977) );
  INVX2 U5070 ( .A(sum[19]), .Y(n5522) );
  INVX2 U5071 ( .A(sum[20]), .Y(n5524) );
  CLKINVXL U5072 ( .A(n6008), .Y(n6016) );
  INVX3 U5073 ( .A(sum[16]), .Y(n5515) );
  INVX2 U5074 ( .A(sum[21]), .Y(n5526) );
  INVX2 U5075 ( .A(sum[10]), .Y(n5501) );
  CLKINVXL U5076 ( .A(n5537), .Y(n5536) );
  OAI2BB1X1 U5077 ( .A0N(n5968), .A1N(n5546), .B0(n5548), .Y(n5969) );
  OAI2BB1X1 U5078 ( .A0N(n5966), .A1N(n5537), .B0(n5540), .Y(n5967) );
  OAI2BB1X1 U5079 ( .A0N(n5965), .A1N(n5532), .B0(n5534), .Y(n5966) );
  OAI2BB1XL U5080 ( .A0N(n5962), .A1N(n5519), .B0(n5522), .Y(n5963) );
  OAI21XL U5081 ( .A0(n5991), .A1(n5990), .B0(n5989), .Y(n5993) );
  CLKINVX2 U5082 ( .A(n6018), .Y(n5994) );
  INVX2 U5083 ( .A(sum[28]), .Y(n5542) );
  INVX1 U5084 ( .A(sum[7]), .Y(n5494) );
  INVX2 U5085 ( .A(sum[12]), .Y(n5506) );
  OAI2BB1XL U5086 ( .A0N(n5960), .A1N(n5510), .B0(n5512), .Y(n5961) );
  OAI2BB1XL U5087 ( .A0N(n5959), .A1N(n5506), .B0(n5508), .Y(n5960) );
  AOI21XL U5088 ( .A0(n5988), .A1(n5987), .B0(n5986), .Y(n5991) );
  CLKINVXL U5089 ( .A(n5985), .Y(n5987) );
  AOI21XL U5090 ( .A0(n5477), .A1(n5480), .B0(n5482), .Y(n2353) );
  INVX2 U5091 ( .A(sum[2]), .Y(n5480) );
  NOR3XL U5092 ( .A(n5974), .B(n5482), .C(n5485), .Y(n5976) );
  OAI2BB1XL U5093 ( .A0N(n6022), .A1N(n6021), .B0(n6020), .Y(n6023) );
  NAND3X1 U5094 ( .A(n6036), .B(n6030), .C(n6029), .Y(n6783) );
  OAI2BB1XL U5095 ( .A0N(N6290), .A1N(n4996), .B0(n6611), .Y(n3468) );
  OAI2BB1XL U5096 ( .A0N(N6249), .A1N(n4995), .B0(n6667), .Y(n3523) );
  OAI2BB1XL U5097 ( .A0N(N6289), .A1N(n4996), .B0(n6612), .Y(n3469) );
  OAI2BB1XL U5098 ( .A0N(N6248), .A1N(n4995), .B0(n6668), .Y(n3524) );
  OAI2BB1XL U5099 ( .A0N(N6372), .A1N(n4999), .B0(n6500), .Y(n3358) );
  OAI2BB1XL U5100 ( .A0N(N6371), .A1N(n4999), .B0(n6501), .Y(n3359) );
  OAI2BB1XL U5101 ( .A0N(N6368), .A1N(n4999), .B0(n6505), .Y(n3362) );
  OAI2BB1XL U5102 ( .A0N(N6208), .A1N(n4994), .B0(n6723), .Y(n3578) );
  OAI2BB1XL U5103 ( .A0N(N6331), .A1N(n4997), .B0(n6555), .Y(n3413) );
  OAI2BB1XL U5104 ( .A0N(N6207), .A1N(n4994), .B0(n6724), .Y(n3579) );
  OAI2BB1XL U5105 ( .A0N(N6330), .A1N(n4997), .B0(n6556), .Y(n3414) );
  OAI2BB1XL U5106 ( .A0N(N6446), .A1N(n4992), .B0(n6404), .Y(n3256) );
  OAI2BB1XL U5107 ( .A0N(N6250), .A1N(n4995), .B0(n6666), .Y(n3522) );
  OAI2BB1XL U5108 ( .A0N(N6449), .A1N(n4992), .B0(n6399), .Y(n3253) );
  OAI2BB1XL U5109 ( .A0N(N6453), .A1N(n4992), .B0(n6394), .Y(n3249) );
  OAI2BB1XL U5110 ( .A0N(N6450), .A1N(n4992), .B0(n6398), .Y(n3252) );
  OAI2BB1XL U5111 ( .A0N(N6209), .A1N(n4994), .B0(n6722), .Y(n3577) );
  OAI2BB1XL U5112 ( .A0N(N6454), .A1N(n4992), .B0(n6393), .Y(n3248) );
  OAI2BB1XL U5113 ( .A0N(N6413), .A1N(n5000), .B0(n6447), .Y(n3303) );
  OAI2BB1XL U5114 ( .A0N(N6409), .A1N(n5000), .B0(n6452), .Y(n3307) );
  OAI2BB1XL U5115 ( .A0N(N6408), .A1N(n5000), .B0(n6453), .Y(n3308) );
  OAI2BB1XL U5116 ( .A0N(N6245), .A1N(n4995), .B0(n6672), .Y(n3527) );
  OAI2BB1XL U5117 ( .A0N(N6445), .A1N(n4992), .B0(n6405), .Y(n3257) );
  OAI2BB1XL U5118 ( .A0N(N6412), .A1N(n5000), .B0(n6448), .Y(n3304) );
  OAI2BB1XL U5119 ( .A0N(N6204), .A1N(n4994), .B0(n6728), .Y(n3582) );
  OAI2BB1XL U5120 ( .A0N(N6455), .A1N(n4992), .B0(n6392), .Y(n3247) );
  OAI2BB1XL U5121 ( .A0N(N6373), .A1N(n4999), .B0(n6499), .Y(n3357) );
  OAI2BB1XL U5122 ( .A0N(N6286), .A1N(n4996), .B0(n6616), .Y(n3472) );
  OAI2BB1XL U5123 ( .A0N(N6490), .A1N(n4993), .B0(n6345), .Y(n3198) );
  OAI2BB1XL U5124 ( .A0N(N6287), .A1N(n4996), .B0(n6615), .Y(n3471) );
  OAI2BB1XL U5125 ( .A0N(N6327), .A1N(n4997), .B0(n6561), .Y(n3417) );
  OAI2BB1XL U5126 ( .A0N(N6405), .A1N(n5000), .B0(n6458), .Y(n3311) );
  OAI2BB1XL U5127 ( .A0N(N6494), .A1N(n4993), .B0(n6340), .Y(n3194) );
  OAI2BB1XL U5128 ( .A0N(N6491), .A1N(n4993), .B0(n6344), .Y(n3197) );
  OAI2BB1XL U5129 ( .A0N(N6451), .A1N(n4992), .B0(n6397), .Y(n3251) );
  OAI2BB1XL U5130 ( .A0N(N6240), .A1N(n4995), .B0(n6679), .Y(n3532) );
  OAI2BB1XL U5131 ( .A0N(N6282), .A1N(n4996), .B0(n6622), .Y(n3476) );
  OAI2BB1XL U5132 ( .A0N(N6323), .A1N(n4997), .B0(n6567), .Y(n3421) );
  OAI2BB1XL U5133 ( .A0N(N6495), .A1N(n4993), .B0(n6339), .Y(n3193) );
  OAI2BB1XL U5134 ( .A0N(N6487), .A1N(n4993), .B0(n6350), .Y(n3201) );
  OAI2BB1XL U5135 ( .A0N(N6241), .A1N(n4995), .B0(n6678), .Y(n3531) );
  OAI2BB1XL U5136 ( .A0N(N6281), .A1N(n4996), .B0(n6623), .Y(n3477) );
  OAI2BB1XL U5137 ( .A0N(N6410), .A1N(n5000), .B0(n6451), .Y(n3306) );
  OAI2BB1XL U5138 ( .A0N(N6486), .A1N(n4993), .B0(n6351), .Y(n3202) );
  OAI2BB1XL U5139 ( .A0N(N6246), .A1N(n4995), .B0(n6671), .Y(n3526) );
  OAI2BB1XL U5140 ( .A0N(N6364), .A1N(n4999), .B0(n6511), .Y(n3366) );
  OAI2BB1XL U5141 ( .A0N(N6404), .A1N(n5000), .B0(n6459), .Y(n3312) );
  OAI2BB1XL U5142 ( .A0N(N6496), .A1N(n4993), .B0(n6338), .Y(n3192) );
  OAI2BB1XL U5143 ( .A0N(N6205), .A1N(n4994), .B0(n6727), .Y(n3581) );
  OAI2BB1XL U5144 ( .A0N(N6414), .A1N(n5000), .B0(n6446), .Y(n3302) );
  OAI2BB1XL U5145 ( .A0N(N6200), .A1N(n4994), .B0(n6734), .Y(n3586) );
  OAI2BB1XL U5146 ( .A0N(N6363), .A1N(n4999), .B0(n6512), .Y(n3367) );
  OAI2BB1XL U5147 ( .A0N(N6322), .A1N(n4997), .B0(n6568), .Y(n3422) );
  OAI2BB1XL U5148 ( .A0N(N6492), .A1N(n4993), .B0(n6343), .Y(n3196) );
  OAI2BB1XL U5149 ( .A0N(N6199), .A1N(n4994), .B0(n6735), .Y(n3587) );
  OAI2BB1XL U5150 ( .A0N(N6237), .A1N(n4995), .B0(n6684), .Y(n3535) );
  OAI2BB1XL U5151 ( .A0N(N6319), .A1N(n4997), .B0(n6572), .Y(n3425) );
  OAI2BB1XL U5152 ( .A0N(N6359), .A1N(n4999), .B0(n6517), .Y(n3371) );
  OAI2BB1XL U5153 ( .A0N(N6196), .A1N(n4994), .B0(n6739), .Y(n3590) );
  OAI2BB1XL U5154 ( .A0N(N6278), .A1N(n4996), .B0(n6628), .Y(n3480) );
  OAI2BB1XL U5155 ( .A0N(N6483), .A1N(n4993), .B0(n6356), .Y(n3205) );
  OAI2BB1XL U5156 ( .A0N(N6401), .A1N(n5000), .B0(n6464), .Y(n3315) );
  OAI2BB1XL U5157 ( .A0N(N6442), .A1N(n4992), .B0(n6410), .Y(n3260) );
  OAI221XL U5158 ( .A0(n6788), .A1(n6039), .B0(n5345), .B1(n6037), .C0(n6786), 
        .Y(n3987) );
  OAI2BB1XL U5159 ( .A0N(N6233), .A1N(n4995), .B0(n6689), .Y(n3539) );
  OAI2BB1XL U5160 ( .A0N(N6274), .A1N(n4996), .B0(n6634), .Y(n3484) );
  OAI2BB1XL U5161 ( .A0N(N6232), .A1N(n4995), .B0(n6690), .Y(n3540) );
  OAI2BB1XL U5162 ( .A0N(N6355), .A1N(n4999), .B0(n6523), .Y(n3375) );
  NAND2BX1 U5163 ( .AN(n6138), .B(y_out_sum5[39]), .Y(n6093) );
  NAND2BX1 U5164 ( .AN(n6286), .B(y_out_sum2[39]), .Y(n6240) );
  NAND2BX1 U5165 ( .AN(n6186), .B(y_out_sum4[39]), .Y(n6141) );
  NAND2BX1 U5166 ( .AN(n6336), .B(y_out_sum1[39]), .Y(n6291) );
  NAND2BX1 U5167 ( .AN(n6235), .B(y_out_sum3[39]), .Y(n6190) );
  NAND2BX1 U5168 ( .AN(n6090), .B(y_out_sum6[39]), .Y(n6045) );
  NAND2BX1 U5169 ( .AN(n5949), .B(y_out_sum0[39]), .Y(n5904) );
  NAND2BX1 U5170 ( .AN(n5949), .B(y_out_sum0[37]), .Y(n5906) );
  NAND2BX1 U5171 ( .AN(n6186), .B(y_out_sum4[37]), .Y(n6143) );
  OAI2BB1XL U5172 ( .A0N(N6333), .A1N(n4997), .B0(n6607), .Y(n3451) );
  NAND2BX1 U5173 ( .AN(n5949), .B(y_out_sum0[36]), .Y(n5907) );
  NAND2BX1 U5174 ( .AN(n5949), .B(y_out_sum0[35]), .Y(n5908) );
  NAND2BX1 U5175 ( .AN(n6186), .B(y_out_sum4[35]), .Y(n6145) );
  NAND2BX1 U5176 ( .AN(n6186), .B(y_out_sum4[36]), .Y(n6144) );
  NAND2BX1 U5177 ( .AN(n6235), .B(y_out_sum3[37]), .Y(n6192) );
  NAND2BX1 U5178 ( .AN(n6336), .B(y_out_sum1[37]), .Y(n6293) );
  NAND2BX1 U5179 ( .AN(n5949), .B(y_out_sum0[32]), .Y(n5911) );
  NAND2BX1 U5180 ( .AN(n5949), .B(y_out_sum0[31]), .Y(n5912) );
  NAND2BX1 U5181 ( .AN(n5949), .B(y_out_sum0[33]), .Y(n5910) );
  NAND2BX1 U5182 ( .AN(n6090), .B(y_out_sum6[37]), .Y(n6047) );
  NAND2BX1 U5183 ( .AN(n5949), .B(y_out_sum0[38]), .Y(n5905) );
  NAND2BX1 U5184 ( .AN(n6138), .B(y_out_sum5[38]), .Y(n6094) );
  NAND2BX1 U5185 ( .AN(n6286), .B(y_out_sum2[38]), .Y(n6241) );
  NAND2BX1 U5186 ( .AN(n6235), .B(y_out_sum3[35]), .Y(n6194) );
  NAND2BX1 U5187 ( .AN(n6186), .B(y_out_sum4[38]), .Y(n6142) );
  NAND2BX1 U5188 ( .AN(n6336), .B(y_out_sum1[36]), .Y(n6294) );
  NAND2BX1 U5189 ( .AN(n6336), .B(y_out_sum1[35]), .Y(n6295) );
  NAND2BX1 U5190 ( .AN(n6090), .B(y_out_sum6[36]), .Y(n6048) );
  NAND2BX1 U5191 ( .AN(n6090), .B(y_out_sum6[35]), .Y(n6049) );
  NAND2BX1 U5192 ( .AN(n6235), .B(y_out_sum3[36]), .Y(n6193) );
  OAI2BB1XL U5193 ( .A0N(N6374), .A1N(n4999), .B0(n6551), .Y(n3396) );
  NAND2BX1 U5194 ( .AN(n6286), .B(y_out_sum2[37]), .Y(n6242) );
  NAND2BX1 U5195 ( .AN(n6138), .B(y_out_sum5[37]), .Y(n6095) );
  NAND2BX1 U5196 ( .AN(n6235), .B(y_out_sum3[38]), .Y(n6191) );
  NAND2BX1 U5197 ( .AN(n6336), .B(y_out_sum1[38]), .Y(n6292) );
  NAND2BX1 U5198 ( .AN(n6286), .B(y_out_sum2[35]), .Y(n6244) );
  NAND2BX1 U5199 ( .AN(n6138), .B(y_out_sum5[35]), .Y(n6097) );
  NAND2BX1 U5200 ( .AN(n6336), .B(y_out_sum1[34]), .Y(n6296) );
  NAND2BX1 U5201 ( .AN(n6336), .B(y_out_sum1[31]), .Y(n6299) );
  NAND2BX1 U5202 ( .AN(n6336), .B(y_out_sum1[32]), .Y(n6298) );
  NAND2BX1 U5203 ( .AN(n6336), .B(y_out_sum1[33]), .Y(n6297) );
  NAND2BX1 U5204 ( .AN(n6138), .B(y_out_sum5[36]), .Y(n6096) );
  NAND2BX1 U5205 ( .AN(n5949), .B(y_out_sum0[34]), .Y(n5909) );
  OAI2BB1XL U5206 ( .A0N(N6251), .A1N(n4995), .B0(n6718), .Y(n3561) );
  NAND2BX1 U5207 ( .AN(n6286), .B(y_out_sum2[36]), .Y(n6243) );
  NAND2BX1 U5208 ( .AN(n6090), .B(y_out_sum6[38]), .Y(n6046) );
  OAI2BB1XL U5209 ( .A0N(N6210), .A1N(n4994), .B0(n6773), .Y(n3616) );
  NAND2BX1 U5210 ( .AN(n6235), .B(y_out_sum3[34]), .Y(n6195) );
  NAND2BX1 U5211 ( .AN(n6235), .B(y_out_sum3[32]), .Y(n6197) );
  NAND2BX1 U5212 ( .AN(n6235), .B(y_out_sum3[31]), .Y(n6198) );
  NAND2BX1 U5213 ( .AN(n6235), .B(y_out_sum3[33]), .Y(n6196) );
  OAI2BB1XL U5214 ( .A0N(N6288), .A1N(n4996), .B0(n6614), .Y(n3470) );
  NAND2BX1 U5215 ( .AN(n6138), .B(y_out_sum5[31]), .Y(n6101) );
  NAND2BX1 U5216 ( .AN(n6138), .B(y_out_sum5[34]), .Y(n6098) );
  NAND2BX1 U5217 ( .AN(n6138), .B(y_out_sum5[33]), .Y(n6099) );
  NAND2BX1 U5218 ( .AN(n6138), .B(y_out_sum5[32]), .Y(n6100) );
  OAI2BB1XL U5219 ( .A0N(N6247), .A1N(n4995), .B0(n6670), .Y(n3525) );
  NAND2BX1 U5220 ( .AN(n5949), .B(y_out_sum0[30]), .Y(n5913) );
  OAI2BB1XL U5221 ( .A0N(N6366), .A1N(n4999), .B0(n6508), .Y(n3364) );
  OAI2BB1XL U5222 ( .A0N(N6370), .A1N(n4999), .B0(n6503), .Y(n3360) );
  NAND2BX1 U5223 ( .AN(n6138), .B(y_out_sum5[29]), .Y(n6103) );
  NAND2BX1 U5224 ( .AN(n6286), .B(y_out_sum2[31]), .Y(n6248) );
  NAND2BX1 U5225 ( .AN(n6286), .B(y_out_sum2[34]), .Y(n6245) );
  NAND2BX1 U5226 ( .AN(n6286), .B(y_out_sum2[32]), .Y(n6247) );
  NAND2BX1 U5227 ( .AN(n6286), .B(y_out_sum2[33]), .Y(n6246) );
  OAI2BB1XL U5228 ( .A0N(N6329), .A1N(n4997), .B0(n6558), .Y(n3415) );
  OAI2BB1XL U5229 ( .A0N(N6206), .A1N(n4994), .B0(n6726), .Y(n3580) );
  OAI2BB1XL U5230 ( .A0N(N6332), .A1N(n4997), .B0(n6554), .Y(n3412) );
  NAND2BX1 U5231 ( .AN(n6186), .B(y_out_sum4[34]), .Y(n6146) );
  NAND2BX1 U5232 ( .AN(n6138), .B(y_out_sum5[28]), .Y(n6104) );
  NAND2BX1 U5233 ( .AN(n6138), .B(y_out_sum5[27]), .Y(n6105) );
  NAND2BX1 U5234 ( .AN(n6138), .B(y_out_sum5[30]), .Y(n6102) );
  NAND2BX1 U5235 ( .AN(n6186), .B(y_out_sum4[31]), .Y(n6149) );
  NAND2BX1 U5236 ( .AN(n6186), .B(y_out_sum4[33]), .Y(n6147) );
  NAND2BX1 U5237 ( .AN(n6186), .B(y_out_sum4[32]), .Y(n6148) );
  OAI2BB1XL U5238 ( .A0N(N6415), .A1N(n5000), .B0(n6497), .Y(n3341) );
  OAI2BB1XL U5239 ( .A0N(N6448), .A1N(n4992), .B0(n6401), .Y(n3254) );
  NAND2BX1 U5240 ( .AN(n5949), .B(y_out_sum0[29]), .Y(n5914) );
  OAI2BB1XL U5241 ( .A0N(N6452), .A1N(n4992), .B0(n6396), .Y(n3250) );
  NAND2BX1 U5242 ( .AN(n6090), .B(y_out_sum6[34]), .Y(n6050) );
  NAND2BX1 U5243 ( .AN(n5949), .B(y_out_sum0[28]), .Y(n5915) );
  NAND2BX1 U5244 ( .AN(n5949), .B(y_out_sum0[27]), .Y(n5916) );
  NAND2BX1 U5245 ( .AN(n6138), .B(y_out_sum5[26]), .Y(n6106) );
  NAND2BX1 U5246 ( .AN(n6090), .B(y_out_sum6[29]), .Y(n6055) );
  OAI2BB1XL U5247 ( .A0N(N6407), .A1N(n5000), .B0(n6455), .Y(n3309) );
  OAI2BB1XL U5248 ( .A0N(N6411), .A1N(n5000), .B0(n6450), .Y(n3305) );
  OAI2BB1XL U5249 ( .A0N(N6243), .A1N(n4995), .B0(n6675), .Y(n3529) );
  NAND2BX1 U5250 ( .AN(n6090), .B(y_out_sum6[31]), .Y(n6053) );
  NAND2BX1 U5251 ( .AN(n6090), .B(y_out_sum6[33]), .Y(n6051) );
  NAND2BX1 U5252 ( .AN(n6090), .B(y_out_sum6[32]), .Y(n6052) );
  OAI2BB1XL U5253 ( .A0N(N6444), .A1N(n4992), .B0(n6407), .Y(n3258) );
  OAI2BB1XL U5254 ( .A0N(N6328), .A1N(n4997), .B0(n6560), .Y(n3416) );
  NAND2BX1 U5255 ( .AN(n6186), .B(y_out_sum4[28]), .Y(n6152) );
  OAI2BB1XL U5256 ( .A0N(N6202), .A1N(n4994), .B0(n6731), .Y(n3584) );
  NAND2BX1 U5257 ( .AN(n6090), .B(y_out_sum6[28]), .Y(n6056) );
  NAND2BX1 U5258 ( .AN(n6090), .B(y_out_sum6[27]), .Y(n6057) );
  NAND2BX1 U5259 ( .AN(n6336), .B(y_out_sum1[30]), .Y(n6300) );
  NAND2BX1 U5260 ( .AN(n6186), .B(y_out_sum4[29]), .Y(n6151) );
  OAI2BB1XL U5261 ( .A0N(N6284), .A1N(n4996), .B0(n6619), .Y(n3474) );
  OAI2BB1XL U5262 ( .A0N(N6489), .A1N(n4993), .B0(n6347), .Y(n3199) );
  OAI2BB1XL U5263 ( .A0N(N6493), .A1N(n4993), .B0(n6342), .Y(n3195) );
  NAND2BX1 U5264 ( .AN(n6186), .B(y_out_sum4[30]), .Y(n6150) );
  OAI2BB1XL U5265 ( .A0N(N6325), .A1N(n4997), .B0(n6564), .Y(n3419) );
  NAND2BX1 U5266 ( .AN(n6235), .B(y_out_sum3[30]), .Y(n6199) );
  NAND2BX1 U5267 ( .AN(n5949), .B(y_out_sum0[26]), .Y(n5917) );
  NAND2BX1 U5268 ( .AN(n6186), .B(y_out_sum4[27]), .Y(n6153) );
  OAI2BB1XL U5269 ( .A0N(N6447), .A1N(n4992), .B0(n6403), .Y(n3255) );
  OAI2BB1XL U5270 ( .A0N(N6280), .A1N(n4996), .B0(n6625), .Y(n3478) );
  OAI2BB1XL U5271 ( .A0N(N6443), .A1N(n4992), .B0(n6409), .Y(n3259) );
  OAI2BB1XL U5272 ( .A0N(N6485), .A1N(n4993), .B0(n6353), .Y(n3203) );
  NAND2BX1 U5273 ( .AN(n6090), .B(y_out_sum6[26]), .Y(n6058) );
  OAI2BB1XL U5274 ( .A0N(N6239), .A1N(n4995), .B0(n6681), .Y(n3533) );
  NAND2BX1 U5275 ( .AN(n6286), .B(y_out_sum2[30]), .Y(n6249) );
  OAI2BB1XL U5276 ( .A0N(N6406), .A1N(n5000), .B0(n6457), .Y(n3310) );
  OAI2BB1XL U5277 ( .A0N(N6242), .A1N(n4995), .B0(n6677), .Y(n3530) );
  OAI2BB1XL U5278 ( .A0N(N6403), .A1N(n5000), .B0(n6461), .Y(n3313) );
  OAI2BB1XL U5279 ( .A0N(N6362), .A1N(n4999), .B0(n6514), .Y(n3368) );
  OAI2BB1XL U5280 ( .A0N(N6201), .A1N(n4994), .B0(n6733), .Y(n3585) );
  OAI2BB1XL U5281 ( .A0N(N6321), .A1N(n4997), .B0(n6570), .Y(n3423) );
  NAND2BX1 U5282 ( .AN(n6186), .B(y_out_sum4[26]), .Y(n6154) );
  OAI2BB1XL U5283 ( .A0N(N6488), .A1N(n4993), .B0(n6349), .Y(n3200) );
  OAI2BB1XL U5284 ( .A0N(N6283), .A1N(n4996), .B0(n6621), .Y(n3475) );
  NAND2BX1 U5285 ( .AN(n6090), .B(y_out_sum6[30]), .Y(n6054) );
  OAI2BB1XL U5286 ( .A0N(N6279), .A1N(n4996), .B0(n6627), .Y(n3479) );
  OAI2BB1XL U5287 ( .A0N(N6324), .A1N(n4997), .B0(n6566), .Y(n3420) );
  OAI2BB1XL U5288 ( .A0N(N6484), .A1N(n4993), .B0(n6355), .Y(n3204) );
  OAI2BB1XL U5289 ( .A0N(N6238), .A1N(n4995), .B0(n6683), .Y(n3534) );
  OAI2BB1XL U5290 ( .A0N(N6198), .A1N(n4994), .B0(n6737), .Y(n3588) );
  OAI2BB1XL U5291 ( .A0N(N6402), .A1N(n5000), .B0(n6463), .Y(n3314) );
  OAI2BB1XL U5292 ( .A0N(N6361), .A1N(n4999), .B0(n6515), .Y(n3369) );
  OAI2BB1XL U5293 ( .A0N(N6320), .A1N(n4997), .B0(n6571), .Y(n3424) );
  NAND2BX1 U5294 ( .AN(n6090), .B(y_out_sum6[24]), .Y(n6060) );
  NAND2BX1 U5295 ( .AN(n6090), .B(y_out_sum6[25]), .Y(n6059) );
  OAI221X1 U5296 ( .A0(n5956), .A1(n6039), .B0(n5346), .B1(n6037), .C0(n6784), 
        .Y(n3989) );
  OAI2BB1XL U5297 ( .A0N(N6197), .A1N(n4994), .B0(n6738), .Y(n3589) );
  NAND2BX1 U5298 ( .AN(n6235), .B(y_out_sum3[27]), .Y(n6202) );
  NAND2BX1 U5299 ( .AN(n6286), .B(y_out_sum2[29]), .Y(n6250) );
  NAND2BX1 U5300 ( .AN(n6235), .B(y_out_sum3[29]), .Y(n6200) );
  NAND2BX1 U5301 ( .AN(n5949), .B(y_out_sum0[24]), .Y(n5919) );
  NAND2BX1 U5302 ( .AN(n5949), .B(y_out_sum0[25]), .Y(n5918) );
  NAND2BX1 U5303 ( .AN(n6235), .B(y_out_sum3[28]), .Y(n6201) );
  NAND2BX1 U5304 ( .AN(n6286), .B(y_out_sum2[28]), .Y(n6251) );
  NAND2BX1 U5305 ( .AN(n6286), .B(y_out_sum2[26]), .Y(n6253) );
  NAND2BX1 U5306 ( .AN(n6336), .B(y_out_sum1[29]), .Y(n6301) );
  NAND2BX1 U5307 ( .AN(n6286), .B(y_out_sum2[27]), .Y(n6252) );
  NAND2BX1 U5308 ( .AN(n6186), .B(y_out_sum4[24]), .Y(n6156) );
  NAND2BX1 U5309 ( .AN(n6286), .B(y_out_sum2[24]), .Y(n6255) );
  NAND2BX1 U5310 ( .AN(n6286), .B(y_out_sum2[25]), .Y(n6254) );
  NAND2BX1 U5311 ( .AN(n6186), .B(y_out_sum4[25]), .Y(n6155) );
  NAND2BX1 U5312 ( .AN(n6138), .B(y_out_sum5[25]), .Y(n6107) );
  NAND2BX1 U5313 ( .AN(n6235), .B(y_out_sum3[24]), .Y(n6205) );
  NAND2BX1 U5314 ( .AN(n6235), .B(y_out_sum3[25]), .Y(n6204) );
  NAND2BX1 U5315 ( .AN(n6336), .B(y_out_sum1[28]), .Y(n6302) );
  NAND2BX1 U5316 ( .AN(n6336), .B(y_out_sum1[27]), .Y(n6303) );
  NAND2BX1 U5317 ( .AN(n6138), .B(y_out_sum5[24]), .Y(n6108) );
  NAND2BX1 U5318 ( .AN(n6235), .B(y_out_sum3[26]), .Y(n6203) );
  NAND2BX1 U5319 ( .AN(n6090), .B(y_out_sum6[23]), .Y(n6061) );
  NAND2BX1 U5320 ( .AN(n6336), .B(y_out_sum1[26]), .Y(n6304) );
  OAI2BB1XL U5321 ( .A0N(n2839), .A1N(n6787), .B0(n6779), .Y(n3176) );
  NAND2BX1 U5322 ( .AN(n5949), .B(y_out_sum0[23]), .Y(n5920) );
  NAND2BX1 U5323 ( .AN(n6336), .B(y_out_sum1[24]), .Y(n6306) );
  NAND2BX1 U5324 ( .AN(n6336), .B(y_out_sum1[25]), .Y(n6305) );
  NAND2BX1 U5325 ( .AN(n6286), .B(y_out_sum2[23]), .Y(n6256) );
  NAND2BX1 U5326 ( .AN(n6186), .B(y_out_sum4[23]), .Y(n6157) );
  NAND2BX1 U5327 ( .AN(n6235), .B(y_out_sum3[23]), .Y(n6206) );
  OAI2BB1XL U5328 ( .A0N(N6235), .A1N(n4995), .B0(n6687), .Y(n3537) );
  NAND2BX1 U5329 ( .AN(n6138), .B(y_out_sum5[23]), .Y(n6109) );
  OAI2BB1XL U5330 ( .A0N(N6317), .A1N(n4997), .B0(n6575), .Y(n3427) );
  OAI2BB1XL U5331 ( .A0N(N6358), .A1N(n4999), .B0(n6519), .Y(n3372) );
  OAI2BB1XL U5332 ( .A0N(N6194), .A1N(n4994), .B0(n6742), .Y(n3592) );
  OAI2BB1XL U5333 ( .A0N(n6787), .A1N(n2841), .B0(n6785), .Y(n3174) );
  OAI2BB1XL U5334 ( .A0N(N6276), .A1N(n4996), .B0(n6631), .Y(n3482) );
  NAND2BX1 U5335 ( .AN(n5949), .B(y_out_sum0[22]), .Y(n5921) );
  NAND2BX1 U5336 ( .AN(n6336), .B(y_out_sum1[23]), .Y(n6307) );
  NAND2BX1 U5337 ( .AN(n6138), .B(y_out_sum5[22]), .Y(n6110) );
  NAND2BX1 U5338 ( .AN(n6286), .B(y_out_sum2[22]), .Y(n6257) );
  NAND2BX1 U5339 ( .AN(n6186), .B(y_out_sum4[22]), .Y(n6158) );
  NAND2BX1 U5340 ( .AN(n6336), .B(y_out_sum1[22]), .Y(n6308) );
  NAND2BX1 U5341 ( .AN(n6090), .B(y_out_sum6[22]), .Y(n6062) );
  NAND2BX1 U5342 ( .AN(n6235), .B(y_out_sum3[22]), .Y(n6207) );
  OAI2BB1XL U5343 ( .A0N(N6234), .A1N(n4995), .B0(n6688), .Y(n3538) );
  OAI2BB1XL U5344 ( .A0N(N6316), .A1N(n4997), .B0(n6577), .Y(n3428) );
  OAI2BB1XL U5345 ( .A0N(n6787), .A1N(n2840), .B0(n6786), .Y(n3175) );
  OAI2BB1XL U5346 ( .A0N(N6357), .A1N(n4999), .B0(n6521), .Y(n3373) );
  OAI2BB1XL U5347 ( .A0N(N6193), .A1N(n4994), .B0(n6743), .Y(n3593) );
  OAI2BB1XL U5348 ( .A0N(N6481), .A1N(n4993), .B0(n6358), .Y(n3207) );
  OAI2BB1XL U5349 ( .A0N(N6399), .A1N(n5000), .B0(n6466), .Y(n3317) );
  NAND2BX1 U5350 ( .AN(n6090), .B(y_out_sum6[21]), .Y(n6063) );
  OAI2BB1XL U5351 ( .A0N(N6440), .A1N(n4992), .B0(n6412), .Y(n3262) );
  NAND2BX1 U5352 ( .AN(n6286), .B(y_out_sum2[21]), .Y(n6258) );
  NAND2BX1 U5353 ( .AN(n6138), .B(y_out_sum5[21]), .Y(n6111) );
  NAND2BX1 U5354 ( .AN(n6186), .B(y_out_sum4[21]), .Y(n6159) );
  OAI2BB1XL U5355 ( .A0N(N6439), .A1N(n4992), .B0(n6413), .Y(n3263) );
  NAND2BX1 U5356 ( .AN(n6235), .B(y_out_sum3[21]), .Y(n6208) );
  NAND2BX1 U5357 ( .AN(n5949), .B(y_out_sum0[21]), .Y(n5922) );
  NAND2BX1 U5358 ( .AN(n6336), .B(y_out_sum1[21]), .Y(n6309) );
  OAI2BB1XL U5359 ( .A0N(N6480), .A1N(n4993), .B0(n6359), .Y(n3208) );
  NAND2BX1 U5360 ( .AN(n6336), .B(y_out_sum1[20]), .Y(n6310) );
  NAND2BX1 U5361 ( .AN(n5949), .B(y_out_sum0[20]), .Y(n5923) );
  OAI2BB1XL U5362 ( .A0N(N6398), .A1N(n5000), .B0(n6467), .Y(n3318) );
  NAND2BX1 U5363 ( .AN(n6138), .B(y_out_sum5[20]), .Y(n6112) );
  NAND2BX1 U5364 ( .AN(n6286), .B(y_out_sum2[20]), .Y(n6259) );
  NAND2BX1 U5365 ( .AN(n6186), .B(y_out_sum4[20]), .Y(n6160) );
  NAND2BX1 U5366 ( .AN(n6090), .B(y_out_sum6[20]), .Y(n6064) );
  NAND2BX1 U5367 ( .AN(n6235), .B(y_out_sum3[20]), .Y(n6209) );
  NAND2BX1 U5368 ( .AN(n5949), .B(y_out_sum0[17]), .Y(n5928) );
  NAND2BX1 U5369 ( .AN(n6605), .B(y_out_sum10[17]), .Y(n6582) );
  NAND2BX1 U5370 ( .AN(n6286), .B(y_out_sum2[17]), .Y(n6264) );
  NAND2BX1 U5371 ( .AN(n6138), .B(y_out_sum5[17]), .Y(n6117) );
  NAND2BX1 U5372 ( .AN(n6235), .B(y_out_sum3[17]), .Y(n6214) );
  NAND2BX1 U5373 ( .AN(n6186), .B(y_out_sum4[17]), .Y(n6165) );
  NAND2BX1 U5374 ( .AN(n6090), .B(y_out_sum6[17]), .Y(n6069) );
  NAND2BX1 U5375 ( .AN(n6661), .B(y_out_sum9[17]), .Y(n6638) );
  NAND2BX1 U5376 ( .AN(n6771), .B(y_out_sum7[17]), .Y(n6748) );
  NAND2BX1 U5377 ( .AN(n6549), .B(y_out_sum11[17]), .Y(n6526) );
  NAND2BX1 U5378 ( .AN(n6716), .B(y_out_sum8[17]), .Y(n6693) );
  NAND2BX1 U5379 ( .AN(n6336), .B(y_out_sum1[17]), .Y(n6315) );
  NAND2BX1 U5380 ( .AN(n6441), .B(y_out_sum13[17]), .Y(n6418) );
  NAND2BX1 U5381 ( .AN(n6387), .B(y_out_sum14[17]), .Y(n6364) );
  NAND2BX1 U5382 ( .AN(n6495), .B(y_out_sum12[17]), .Y(n6472) );
  NAND2BX1 U5383 ( .AN(n6138), .B(y_out_sum5[14]), .Y(n6122) );
  NAND2BX1 U5384 ( .AN(n6186), .B(y_out_sum4[14]), .Y(n6170) );
  NAND2BX1 U5385 ( .AN(n6090), .B(y_out_sum6[14]), .Y(n6074) );
  NAND2BX1 U5386 ( .AN(n6235), .B(y_out_sum3[14]), .Y(n6219) );
  NAND2BX1 U5387 ( .AN(n5949), .B(y_out_sum0[14]), .Y(n5933) );
  NAND2BX1 U5388 ( .AN(n6336), .B(y_out_sum1[14]), .Y(n6320) );
  NAND2BX1 U5389 ( .AN(n6286), .B(y_out_sum2[14]), .Y(n6269) );
  NAND2BX1 U5390 ( .AN(n6138), .B(y_out_sum5[13]), .Y(n6123) );
  NAND2BX1 U5391 ( .AN(n6387), .B(y_out_sum14[13]), .Y(n6369) );
  NAND2BX1 U5392 ( .AN(n6090), .B(y_out_sum6[13]), .Y(n6075) );
  NAND2BX1 U5393 ( .AN(n6186), .B(y_out_sum4[13]), .Y(n6171) );
  NAND2BX1 U5394 ( .AN(n6716), .B(y_out_sum8[13]), .Y(n6698) );
  NAND2BX1 U5395 ( .AN(n6661), .B(y_out_sum9[13]), .Y(n6643) );
  NAND2BX1 U5396 ( .AN(n6771), .B(y_out_sum7[13]), .Y(n6753) );
  NAND2BX1 U5397 ( .AN(n6549), .B(y_out_sum11[13]), .Y(n6531) );
  NAND2BX1 U5398 ( .AN(n6495), .B(y_out_sum12[13]), .Y(n6477) );
  NAND2BX1 U5399 ( .AN(n6605), .B(y_out_sum10[13]), .Y(n6587) );
  NAND2BX1 U5400 ( .AN(n6441), .B(y_out_sum13[13]), .Y(n6423) );
  NAND2BX1 U5401 ( .AN(n5949), .B(y_out_sum0[13]), .Y(n5934) );
  NAND2BX1 U5402 ( .AN(n6235), .B(y_out_sum3[13]), .Y(n6220) );
  NAND2BX1 U5403 ( .AN(n6286), .B(y_out_sum2[13]), .Y(n6270) );
  NAND2BX1 U5404 ( .AN(n6336), .B(y_out_sum1[13]), .Y(n6321) );
  NAND2BX1 U5405 ( .AN(n6138), .B(y_out_sum5[12]), .Y(n6124) );
  NAND2BX1 U5406 ( .AN(n6387), .B(y_out_sum14[12]), .Y(n6370) );
  NAND2BX1 U5407 ( .AN(n6441), .B(y_out_sum13[12]), .Y(n6424) );
  NAND2BX1 U5408 ( .AN(n6186), .B(y_out_sum4[12]), .Y(n6172) );
  NAND2BX1 U5409 ( .AN(n6090), .B(y_out_sum6[12]), .Y(n6076) );
  NAND2BX1 U5410 ( .AN(n6661), .B(y_out_sum9[12]), .Y(n6644) );
  NAND2BX1 U5411 ( .AN(n6771), .B(y_out_sum7[12]), .Y(n6754) );
  NAND2BX1 U5412 ( .AN(n6549), .B(y_out_sum11[12]), .Y(n6532) );
  NAND2BX1 U5413 ( .AN(n6495), .B(y_out_sum12[12]), .Y(n6478) );
  NAND2BX1 U5414 ( .AN(n6716), .B(y_out_sum8[12]), .Y(n6699) );
  NAND2BX1 U5415 ( .AN(n6605), .B(y_out_sum10[12]), .Y(n6588) );
  NAND2BX1 U5416 ( .AN(n5949), .B(y_out_sum0[12]), .Y(n5935) );
  NAND2BX1 U5417 ( .AN(n6286), .B(y_out_sum2[12]), .Y(n6271) );
  NAND2BX1 U5418 ( .AN(n6138), .B(y_out_sum5[11]), .Y(n6125) );
  NAND2BX1 U5419 ( .AN(n6336), .B(y_out_sum1[12]), .Y(n6322) );
  NAND2BX1 U5420 ( .AN(n6235), .B(y_out_sum3[12]), .Y(n6221) );
  NAND2BX1 U5421 ( .AN(n6186), .B(y_out_sum4[11]), .Y(n6173) );
  NAND2BX1 U5422 ( .AN(n6090), .B(y_out_sum6[11]), .Y(n6077) );
  NAND2BX1 U5423 ( .AN(n5949), .B(y_out_sum0[11]), .Y(n5936) );
  NAND2BX1 U5424 ( .AN(n6286), .B(y_out_sum2[11]), .Y(n6272) );
  NAND2BX1 U5425 ( .AN(n6235), .B(y_out_sum3[11]), .Y(n6222) );
  NAND2BX1 U5426 ( .AN(n6138), .B(y_out_sum5[10]), .Y(n6126) );
  NAND2BX1 U5427 ( .AN(n6336), .B(y_out_sum1[11]), .Y(n6323) );
  NAND2BX1 U5428 ( .AN(n6186), .B(y_out_sum4[10]), .Y(n6174) );
  NAND2BX1 U5429 ( .AN(n6090), .B(y_out_sum6[10]), .Y(n6078) );
  NAND2BX1 U5430 ( .AN(n5949), .B(y_out_sum0[10]), .Y(n5937) );
  NAND2BX1 U5431 ( .AN(n6186), .B(y_out_sum4[9]), .Y(n6175) );
  NAND2BX1 U5432 ( .AN(n6090), .B(y_out_sum6[9]), .Y(n6079) );
  NAND2BX1 U5433 ( .AN(n6661), .B(y_out_sum9[9]), .Y(n6647) );
  NAND2BX1 U5434 ( .AN(n6771), .B(y_out_sum7[9]), .Y(n6757) );
  NAND2BX1 U5435 ( .AN(n6549), .B(y_out_sum11[9]), .Y(n6535) );
  NAND2BX1 U5436 ( .AN(n6495), .B(y_out_sum12[9]), .Y(n6481) );
  NAND2BX1 U5437 ( .AN(n6716), .B(y_out_sum8[9]), .Y(n6702) );
  NAND2BX1 U5438 ( .AN(n6605), .B(y_out_sum10[9]), .Y(n6591) );
  NAND2BX1 U5439 ( .AN(n6441), .B(y_out_sum13[9]), .Y(n6427) );
  NAND2BX1 U5440 ( .AN(n6387), .B(y_out_sum14[9]), .Y(n6373) );
  NAND2BX1 U5441 ( .AN(n5949), .B(y_out_sum0[9]), .Y(n5938) );
  NAND2BX1 U5442 ( .AN(n6138), .B(y_out_sum5[9]), .Y(n6127) );
  NAND2BX1 U5443 ( .AN(n6336), .B(y_out_sum1[10]), .Y(n6324) );
  NAND2BX1 U5444 ( .AN(n6286), .B(y_out_sum2[10]), .Y(n6273) );
  NAND2BX1 U5445 ( .AN(n6235), .B(y_out_sum3[10]), .Y(n6223) );
  NAND2BX1 U5446 ( .AN(n6186), .B(y_out_sum4[8]), .Y(n6176) );
  NAND2BX1 U5447 ( .AN(n6138), .B(y_out_sum5[8]), .Y(n6128) );
  NAND2BX1 U5448 ( .AN(n6090), .B(y_out_sum6[8]), .Y(n6080) );
  NAND2BX1 U5449 ( .AN(n6661), .B(y_out_sum9[8]), .Y(n6648) );
  NAND2BX1 U5450 ( .AN(n6771), .B(y_out_sum7[8]), .Y(n6758) );
  NAND2BX1 U5451 ( .AN(n6549), .B(y_out_sum11[8]), .Y(n6536) );
  NAND2BX1 U5452 ( .AN(n6495), .B(y_out_sum12[8]), .Y(n6482) );
  NAND2BX1 U5453 ( .AN(n6605), .B(y_out_sum10[8]), .Y(n6592) );
  NAND2BX1 U5454 ( .AN(n6441), .B(y_out_sum13[8]), .Y(n6428) );
  NAND2BX1 U5455 ( .AN(n6387), .B(y_out_sum14[8]), .Y(n6374) );
  NAND2BX1 U5456 ( .AN(n6716), .B(y_out_sum8[8]), .Y(n6703) );
  NAND2BX1 U5457 ( .AN(n5949), .B(y_out_sum0[8]), .Y(n5939) );
  NAND2BX1 U5458 ( .AN(n6336), .B(y_out_sum1[9]), .Y(n6325) );
  NAND2BX1 U5459 ( .AN(n6286), .B(y_out_sum2[9]), .Y(n6274) );
  NAND2BX1 U5460 ( .AN(n6235), .B(y_out_sum3[9]), .Y(n6224) );
  NAND2BX1 U5461 ( .AN(n6336), .B(y_out_sum1[8]), .Y(n6326) );
  NAND2BX1 U5462 ( .AN(n6286), .B(y_out_sum2[8]), .Y(n6275) );
  NAND2BX1 U5463 ( .AN(n6235), .B(y_out_sum3[8]), .Y(n6225) );
  NAND2BX1 U5464 ( .AN(n6186), .B(y_out_sum4[7]), .Y(n6177) );
  NAND2BX1 U5465 ( .AN(n6138), .B(y_out_sum5[7]), .Y(n6129) );
  NAND2BX1 U5466 ( .AN(n6090), .B(y_out_sum6[7]), .Y(n6081) );
  NAND2BX1 U5467 ( .AN(n5949), .B(y_out_sum0[7]), .Y(n5940) );
  NAND2BX1 U5468 ( .AN(n6186), .B(y_out_sum4[6]), .Y(n6178) );
  NAND2BX1 U5469 ( .AN(n6138), .B(y_out_sum5[6]), .Y(n6130) );
  NAND2BX1 U5470 ( .AN(n6090), .B(y_out_sum6[6]), .Y(n6082) );
  NAND2BX1 U5471 ( .AN(n5949), .B(y_out_sum0[6]), .Y(n5941) );
  NAND2BX1 U5472 ( .AN(n6286), .B(y_out_sum2[7]), .Y(n6276) );
  NAND2BX1 U5473 ( .AN(n6235), .B(y_out_sum3[7]), .Y(n6226) );
  NAND2BX1 U5474 ( .AN(n6336), .B(y_out_sum1[7]), .Y(n6327) );
  NAND2BX1 U5475 ( .AN(n6336), .B(y_out_sum1[6]), .Y(n6328) );
  NAND2BX1 U5476 ( .AN(n6235), .B(y_out_sum3[6]), .Y(n6227) );
  NAND2BX1 U5477 ( .AN(n6286), .B(y_out_sum2[6]), .Y(n6277) );
  NAND2BX1 U5478 ( .AN(n6090), .B(y_out_sum6[5]), .Y(n6083) );
  NAND2BX1 U5479 ( .AN(n6186), .B(y_out_sum4[5]), .Y(n6179) );
  NAND2BX1 U5480 ( .AN(n5949), .B(y_out_sum0[5]), .Y(n5942) );
  NAND2BX1 U5481 ( .AN(n6138), .B(y_out_sum5[5]), .Y(n6131) );
  NAND2BX1 U5482 ( .AN(n6336), .B(y_out_sum1[5]), .Y(n6329) );
  NAND2BX1 U5483 ( .AN(n6286), .B(y_out_sum2[5]), .Y(n6278) );
  NAND2BX1 U5484 ( .AN(n6235), .B(y_out_sum3[5]), .Y(n6228) );
  NAND2BX1 U5485 ( .AN(n6090), .B(y_out_sum6[4]), .Y(n6084) );
  NAND2BX1 U5486 ( .AN(n5949), .B(y_out_sum0[4]), .Y(n5943) );
  NAND2BX1 U5487 ( .AN(n6186), .B(y_out_sum4[4]), .Y(n6180) );
  NAND2BX1 U5488 ( .AN(n6138), .B(y_out_sum5[4]), .Y(n6132) );
  NAND2BX1 U5489 ( .AN(n6286), .B(y_out_sum2[4]), .Y(n6279) );
  NAND2BX1 U5490 ( .AN(n6235), .B(y_out_sum3[4]), .Y(n6229) );
  NAND2BX1 U5491 ( .AN(n6336), .B(y_out_sum1[4]), .Y(n6330) );
  NAND2BX1 U5492 ( .AN(n6286), .B(y_out_sum2[3]), .Y(n6280) );
  NAND2BX1 U5493 ( .AN(n6235), .B(y_out_sum3[3]), .Y(n6230) );
  NAND2BX1 U5494 ( .AN(n6336), .B(y_out_sum1[3]), .Y(n6331) );
  NAND2BX1 U5495 ( .AN(n6186), .B(y_out_sum4[3]), .Y(n6181) );
  NAND2BX1 U5496 ( .AN(n6090), .B(y_out_sum6[3]), .Y(n6085) );
  NAND2BX1 U5497 ( .AN(n5949), .B(y_out_sum0[3]), .Y(n5944) );
  NAND2BX1 U5498 ( .AN(n6138), .B(y_out_sum5[3]), .Y(n6133) );
  NAND2BX1 U5499 ( .AN(n6336), .B(y_out_sum1[2]), .Y(n6332) );
  NAND2BX1 U5500 ( .AN(n6186), .B(y_out_sum4[2]), .Y(n6182) );
  NAND2BX1 U5501 ( .AN(n6138), .B(y_out_sum5[2]), .Y(n6134) );
  NAND2BX1 U5502 ( .AN(n6090), .B(y_out_sum6[2]), .Y(n6086) );
  NAND2BX1 U5503 ( .AN(n6235), .B(y_out_sum3[2]), .Y(n6231) );
  NAND2BX1 U5504 ( .AN(n5949), .B(y_out_sum0[2]), .Y(n5945) );
  NAND2BXL U5505 ( .AN(n5401), .B(x_in5[4]), .Y(n5835) );
  NAND2BXL U5506 ( .AN(n5401), .B(x_in3[13]), .Y(n5876) );
  NAND2BXL U5507 ( .AN(n5401), .B(x_in4[12]), .Y(n5859) );
  NAND2BXL U5508 ( .AN(n5401), .B(x_in4[6]), .Y(n5853) );
  NAND2BXL U5509 ( .AN(n5401), .B(x_in4[9]), .Y(n5856) );
  NAND2BXL U5510 ( .AN(n5401), .B(x_in4[3]), .Y(n5850) );
  NAND2BXL U5511 ( .AN(n5401), .B(x_in4[5]), .Y(n5852) );
  NAND2BXL U5512 ( .AN(n5401), .B(x_in4[7]), .Y(n5854) );
  NAND2BXL U5513 ( .AN(n5401), .B(x_in6[11]), .Y(n5826) );
  NAND2BXL U5514 ( .AN(n5401), .B(x_in6[12]), .Y(n5827) );
  NAND2BXL U5515 ( .AN(n5401), .B(x_in6[13]), .Y(n5828) );
  NAND2BXL U5516 ( .AN(n5401), .B(x_in6[14]), .Y(n5829) );
  NAND2BXL U5517 ( .AN(n5401), .B(x_in6[15]), .Y(n5830) );
  NAND2BXL U5518 ( .AN(n5401), .B(x_in5[10]), .Y(n5841) );
  NAND2BXL U5519 ( .AN(n5401), .B(x_in5[13]), .Y(n5844) );
  NAND2BXL U5520 ( .AN(n5401), .B(x_in5[1]), .Y(n5832) );
  NAND2BXL U5521 ( .AN(n5401), .B(x_in5[2]), .Y(n5833) );
  NAND2BXL U5522 ( .AN(n5401), .B(x_in5[7]), .Y(n5838) );
  NAND2BXL U5523 ( .AN(n5401), .B(x_in5[9]), .Y(n5840) );
  NAND2BXL U5524 ( .AN(n5401), .B(x_in4[10]), .Y(n5857) );
  NAND2BXL U5525 ( .AN(n5401), .B(x_in4[11]), .Y(n5858) );
  NAND2BXL U5526 ( .AN(n5401), .B(x_in4[13]), .Y(n5860) );
  NAND2BXL U5527 ( .AN(n5401), .B(x_in4[14]), .Y(n5861) );
  NAND2BXL U5528 ( .AN(n5401), .B(x_in4[1]), .Y(n5848) );
  NAND2BXL U5529 ( .AN(n5401), .B(x_in4[2]), .Y(n5849) );
  NAND2BXL U5530 ( .AN(n5401), .B(x_in4[4]), .Y(n5851) );
  NAND2BXL U5531 ( .AN(n5401), .B(x_in4[8]), .Y(n5855) );
  NAND2BXL U5532 ( .AN(n5401), .B(x_in5[11]), .Y(n5842) );
  NAND2BXL U5533 ( .AN(n5401), .B(x_in5[12]), .Y(n5843) );
  NAND2BXL U5534 ( .AN(n5401), .B(x_in5[14]), .Y(n5845) );
  NAND2BXL U5535 ( .AN(n5401), .B(x_in5[15]), .Y(n5846) );
  NAND2BXL U5536 ( .AN(n5401), .B(x_in5[3]), .Y(n5834) );
  NAND2BXL U5537 ( .AN(n5401), .B(x_in5[5]), .Y(n5836) );
  NAND2BXL U5538 ( .AN(n5401), .B(x_in5[6]), .Y(n5837) );
  NAND2BXL U5539 ( .AN(n5401), .B(x_in5[8]), .Y(n5839) );
  NAND2BXL U5540 ( .AN(n5400), .B(x_in2[10]), .Y(n5889) );
  NAND2BXL U5541 ( .AN(n5400), .B(x_in2[11]), .Y(n5890) );
  NAND2BXL U5542 ( .AN(n5400), .B(x_in2[12]), .Y(n5891) );
  NAND2BXL U5543 ( .AN(n5400), .B(x_in2[13]), .Y(n5892) );
  NAND2BXL U5544 ( .AN(n5400), .B(x_in2[14]), .Y(n5893) );
  NAND2BXL U5545 ( .AN(n5400), .B(x_in2[15]), .Y(n5894) );
  NAND2BXL U5546 ( .AN(n5400), .B(x_in2[1]), .Y(n5880) );
  NAND2BXL U5547 ( .AN(n5400), .B(x_in2[2]), .Y(n5881) );
  NAND2BXL U5548 ( .AN(n5400), .B(x_in2[3]), .Y(n5882) );
  NAND2BXL U5549 ( .AN(n5400), .B(x_in2[4]), .Y(n5883) );
  NAND2BXL U5550 ( .AN(n5400), .B(x_in2[5]), .Y(n5884) );
  NAND2BXL U5551 ( .AN(n5400), .B(x_in2[6]), .Y(n5885) );
  NAND2BXL U5552 ( .AN(n5400), .B(x_in2[7]), .Y(n5886) );
  NAND2BXL U5553 ( .AN(n5400), .B(x_in2[8]), .Y(n5887) );
  NAND2BXL U5554 ( .AN(n5400), .B(x_in2[9]), .Y(n5888) );
  NAND2BXL U5555 ( .AN(n5400), .B(x_in3[10]), .Y(n5873) );
  NAND2BXL U5556 ( .AN(n5400), .B(x_in3[11]), .Y(n5874) );
  NAND2BXL U5557 ( .AN(n5400), .B(x_in3[12]), .Y(n5875) );
  NAND2BXL U5558 ( .AN(n5400), .B(x_in3[14]), .Y(n5877) );
  NAND2BXL U5559 ( .AN(n5400), .B(x_in3[15]), .Y(n5878) );
  NAND2BXL U5560 ( .AN(n5400), .B(x_in3[1]), .Y(n5864) );
  NAND2BXL U5561 ( .AN(n5400), .B(x_in3[2]), .Y(n5865) );
  NAND2BXL U5562 ( .AN(n5400), .B(x_in3[3]), .Y(n5866) );
  NAND2BXL U5563 ( .AN(n5400), .B(x_in3[4]), .Y(n5867) );
  NAND2BXL U5564 ( .AN(n5400), .B(x_in3[5]), .Y(n5868) );
  NAND2BXL U5565 ( .AN(n5400), .B(x_in3[6]), .Y(n5869) );
  NAND2BXL U5566 ( .AN(n5400), .B(x_in3[7]), .Y(n5870) );
  NAND2BXL U5567 ( .AN(n5400), .B(x_in3[8]), .Y(n5871) );
  NAND2BXL U5568 ( .AN(n5400), .B(x_in3[9]), .Y(n5872) );
  NAND2BXL U5569 ( .AN(n5400), .B(x_in4[15]), .Y(n5862) );
  NAND2BXL U5570 ( .AN(n5401), .B(x_in7[2]), .Y(n5801) );
  NAND2BXL U5571 ( .AN(n5401), .B(x_in6[10]), .Y(n5825) );
  NAND2BXL U5572 ( .AN(n5401), .B(x_in6[1]), .Y(n5816) );
  NAND2BXL U5573 ( .AN(n5401), .B(x_in6[2]), .Y(n5817) );
  NAND2BXL U5574 ( .AN(n5401), .B(x_in6[3]), .Y(n5818) );
  NAND2BXL U5575 ( .AN(n5401), .B(x_in6[4]), .Y(n5819) );
  NAND2BXL U5576 ( .AN(n5401), .B(x_in6[5]), .Y(n5820) );
  NAND2BXL U5577 ( .AN(n5401), .B(x_in6[6]), .Y(n5821) );
  NAND2BXL U5578 ( .AN(n5401), .B(x_in6[7]), .Y(n5822) );
  NAND2BXL U5579 ( .AN(n5401), .B(x_in6[8]), .Y(n5823) );
  NAND2BXL U5580 ( .AN(n5401), .B(x_in6[9]), .Y(n5824) );
  NAND2BXL U5581 ( .AN(n5401), .B(x_in7[10]), .Y(n5809) );
  NAND2BXL U5582 ( .AN(n5396), .B(x_in7[11]), .Y(n5810) );
  NAND2BXL U5583 ( .AN(n5401), .B(x_in7[12]), .Y(n5811) );
  NAND2BXL U5584 ( .AN(n5401), .B(x_in7[13]), .Y(n5812) );
  NAND2BXL U5585 ( .AN(n5401), .B(x_in7[14]), .Y(n5813) );
  NAND2BXL U5586 ( .AN(n5401), .B(x_in7[15]), .Y(n5814) );
  NAND2BXL U5587 ( .AN(n5398), .B(x_in7[1]), .Y(n5800) );
  NAND2BXL U5588 ( .AN(n5398), .B(x_in7[3]), .Y(n5802) );
  NAND2BXL U5589 ( .AN(n5401), .B(x_in7[4]), .Y(n5803) );
  NAND2BXL U5590 ( .AN(n5401), .B(x_in7[5]), .Y(n5804) );
  NAND2BXL U5591 ( .AN(n5396), .B(x_in7[6]), .Y(n5805) );
  NAND2BXL U5592 ( .AN(n5396), .B(x_in7[7]), .Y(n5806) );
  NAND2BXL U5593 ( .AN(n5398), .B(x_in7[8]), .Y(n5807) );
  NAND2BXL U5594 ( .AN(n5398), .B(x_in7[9]), .Y(n5808) );
  OR2X1 U5595 ( .A(n6011), .B(n6008), .Y(n6027) );
  OR2X1 U5596 ( .A(n5986), .B(n5990), .Y(n6008) );
  OR2X1 U5597 ( .A(n5523), .B(n5521), .Y(n5986) );
  OR2X1 U5598 ( .A(n5981), .B(n5985), .Y(n6011) );
  INVX2 U5599 ( .A(n6009), .Y(n6014) );
  INVX2 U5600 ( .A(n5981), .Y(n5982) );
  INVX2 U5601 ( .A(n5977), .Y(n5979) );
  INVX2 U5602 ( .A(n5557), .Y(n5556) );
  OR3X2 U5603 ( .A(n6018), .B(n6007), .C(n5531), .Y(n6028) );
  INVX2 U5604 ( .A(n5517), .Y(n5516) );
  OR2X1 U5605 ( .A(n5527), .B(sum[21]), .Y(n5990) );
  OR2X1 U5606 ( .A(n5978), .B(n5984), .Y(n6009) );
  CLKINVXL U5607 ( .A(n5995), .Y(n5996) );
  OR2X1 U5608 ( .A(n5541), .B(n5539), .Y(n5992) );
  OR2X1 U5609 ( .A(n4973), .B(n5543), .Y(n5998) );
  INVX2 U5610 ( .A(n5526), .Y(n5525) );
  INVX2 U5611 ( .A(n5501), .Y(n5500) );
  INVX2 U5612 ( .A(n5515), .Y(n5514) );
  INVX2 U5613 ( .A(n5501), .Y(n5499) );
  OR2X1 U5614 ( .A(n5536), .B(sum[25]), .Y(n6018) );
  AND2X1 U5615 ( .A(n6016), .B(n6015), .Y(n6017) );
  OAI2BB1X1 U5616 ( .A0N(n6014), .A1N(n6013), .B0(n6012), .Y(n6015) );
  OR2X1 U5617 ( .A(sum[14]), .B(n5507), .Y(n5984) );
  NOR2X1 U5618 ( .A(n5495), .B(n5493), .Y(n4987) );
  INVX2 U5619 ( .A(n5542), .Y(n5541) );
  CLKINVX8 U5620 ( .A(n5544), .Y(n5543) );
  INVX2 U5621 ( .A(n5540), .Y(n5539) );
  INVX2 U5622 ( .A(n5486), .Y(n5484) );
  INVX2 U5623 ( .A(n5506), .Y(n5504) );
  INVX2 U5624 ( .A(n5486), .Y(n5485) );
  INVX2 U5625 ( .A(n5494), .Y(n5493) );
  INVX2 U5626 ( .A(n5506), .Y(n5505) );
  INVX2 U5627 ( .A(n5488), .Y(n5487) );
  INVX2 U5628 ( .A(n5508), .Y(n5507) );
  INVX2 U5629 ( .A(n5491), .Y(n5490) );
  OAI2BB1XL U5630 ( .A0N(n5964), .A1N(n5528), .B0(n5530), .Y(n5965) );
  OAI2BB1X1 U5631 ( .A0N(n5963), .A1N(n5524), .B0(n5526), .Y(n5964) );
  OAI2BB1X1 U5632 ( .A0N(n5961), .A1N(n5515), .B0(n5517), .Y(n5962) );
  OAI2BB1XL U5633 ( .A0N(n5967), .A1N(n5542), .B0(n5544), .Y(n5968) );
  AOI21XL U5634 ( .A0(n5994), .A1(n5993), .B0(n5992), .Y(n5997) );
  NOR2X1 U5635 ( .A(n4977), .B(n5531), .Y(n5989) );
  NAND4XL U5636 ( .A(n4987), .B(n5498), .C(n6010), .D(n5501), .Y(n6013) );
  INVX2 U5637 ( .A(n5480), .Y(n5479) );
  INVX2 U5638 ( .A(sum[26]), .Y(n5537) );
  OAI21XL U5639 ( .A0(n2350), .A1(n5500), .B0(n5503), .Y(n5959) );
  AOI2BB1X1 U5640 ( .A0N(n5495), .A1N(n2351), .B0(sum[9]), .Y(n2350) );
  OAI21X1 U5641 ( .A0(n5984), .A1(n5983), .B0(n5982), .Y(n5988) );
  AOI21X1 U5642 ( .A0(n5980), .A1(n5979), .B0(n5978), .Y(n5983) );
  OAI21X1 U5643 ( .A0(n5976), .A1(n5975), .B0(n4987), .Y(n5980) );
  NAND2XL U5644 ( .A(n5488), .B(n5491), .Y(n5975) );
  NOR2X1 U5645 ( .A(n5477), .B(sum[2]), .Y(n5974) );
  INVX2 U5646 ( .A(n5478), .Y(n5476) );
  CLKINVXL U5647 ( .A(n5478), .Y(n5477) );
  INVX2 U5648 ( .A(n5475), .Y(n5474) );
  INVX2 U5649 ( .A(sum[0]), .Y(n5475) );
  INVX2 U5650 ( .A(n1993), .Y(n7317) );
  OAI2BB1X1 U5651 ( .A0N(n5972), .A1N(n5557), .B0(n4988), .Y(n6779) );
  OAI2BB1X1 U5652 ( .A0N(n5970), .A1N(n5554), .B0(n5566), .Y(n5971) );
  OAI2BB1X1 U5653 ( .A0N(n6024), .A1N(n6023), .B0(n4988), .Y(n6785) );
  CLKINVXL U5654 ( .A(n6006), .Y(n6024) );
  CLKINVXL U5655 ( .A(n6007), .Y(n6022) );
  OAI21XL U5656 ( .A0(n6004), .A1(n6003), .B0(n4988), .Y(n6786) );
  AOI21XL U5657 ( .A0(n6002), .A1(n6001), .B0(n6000), .Y(n6003) );
  CLKINVXL U5658 ( .A(n5999), .Y(n6001) );
  OAI21XL U5659 ( .A0(n5998), .A1(n5997), .B0(n5996), .Y(n6002) );
  INVX2 U5660 ( .A(n5459), .Y(n5442) );
  INVX2 U5661 ( .A(n2777), .Y(n7233) );
  NAND2X1 U5662 ( .A(n7324), .B(n7045), .Y(n1993) );
  INVX2 U5663 ( .A(n1774), .Y(n7219) );
  INVX2 U5664 ( .A(n1859), .Y(n7196) );
  INVX2 U5665 ( .A(n1457), .Y(n7226) );
  INVX2 U5666 ( .A(n2276), .Y(n7210) );
  INVX2 U5667 ( .A(n1404), .Y(n7227) );
  INVX2 U5668 ( .A(n2023), .Y(n7215) );
  INVX2 U5669 ( .A(n1558), .Y(n7224) );
  INVX2 U5670 ( .A(n1714), .Y(n7221) );
  INVX2 U5671 ( .A(n1662), .Y(n7222) );
  INVX2 U5672 ( .A(n1609), .Y(n7223) );
  INVX2 U5673 ( .A(n1509), .Y(n7225) );
  INVX2 U5674 ( .A(n2102), .Y(n7212) );
  INVX2 U5675 ( .A(n1351), .Y(n7228) );
  INVX2 U5676 ( .A(n1941), .Y(n7217) );
  INVX2 U5677 ( .A(n6549), .Y(n5391) );
  INVX2 U5678 ( .A(n2108), .Y(n7321) );
  INVX2 U5679 ( .A(n2686), .Y(n7231) );
  INVX2 U5680 ( .A(n2601), .Y(n7208) );
  INVX2 U5681 ( .A(n5457), .Y(n5441) );
  INVX2 U5682 ( .A(n5458), .Y(n5438) );
  INVX2 U5683 ( .A(n5458), .Y(n5439) );
  INVX2 U5684 ( .A(n5458), .Y(n5437) );
  INVX2 U5685 ( .A(n5459), .Y(n5440) );
  OR2X1 U5686 ( .A(n6036), .B(n6035), .Y(n6782) );
  NOR2X1 U5687 ( .A(sum[39]), .B(n6035), .Y(n4988) );
  INVX2 U5688 ( .A(n2634), .Y(n7174) );
  INVX2 U5689 ( .A(n2723), .Y(n7019) );
  INVX2 U5690 ( .A(n1864), .Y(n7013) );
  AND3X2 U5691 ( .A(n2684), .B(n2681), .C(n2682), .Y(n2556) );
  NOR2BX1 U5692 ( .AN(n2681), .B(n2684), .Y(n2557) );
  INVX2 U5693 ( .A(n2461), .Y(n7045) );
  NOR2X1 U5694 ( .A(n2649), .B(n2650), .Y(n2558) );
  NOR2BX1 U5695 ( .AN(n2647), .B(n2648), .Y(n2559) );
  NAND2X1 U5696 ( .A(n7323), .B(n1863), .Y(n2721) );
  INVX2 U5697 ( .A(n2710), .Y(n7323) );
  INVX2 U5698 ( .A(n1863), .Y(n7324) );
  NAND2X1 U5699 ( .A(n7326), .B(n7025), .Y(n2108) );
  OR2X1 U5700 ( .A(n2580), .B(n7233), .Y(n2591) );
  INVX2 U5701 ( .A(n5431), .Y(n5459) );
  NOR2X1 U5702 ( .A(n1863), .B(n2697), .Y(n1907) );
  NAND2X1 U5703 ( .A(n7034), .B(n2690), .Y(n2666) );
  OAI21X1 U5704 ( .A0(n7025), .A1(n2153), .B0(n6288), .Y(n2690) );
  INVX2 U5705 ( .A(n6288), .Y(n7018) );
  INVX2 U5706 ( .A(n1290), .Y(n7181) );
  NAND3X1 U5707 ( .A(n7019), .B(n7027), .C(n7030), .Y(n2686) );
  INVX2 U5708 ( .A(n2697), .Y(n7043) );
  INVX2 U5709 ( .A(n1301), .Y(n7179) );
  NAND3X1 U5710 ( .A(n7019), .B(n7027), .C(n7029), .Y(n2777) );
  INVX2 U5711 ( .A(n5423), .Y(n5422) );
  INVX2 U5712 ( .A(n5424), .Y(n5421) );
  INVX2 U5713 ( .A(n5424), .Y(n5420) );
  INVX2 U5714 ( .A(n5424), .Y(n5419) );
  INVX2 U5715 ( .A(n5423), .Y(n5418) );
  INVX2 U5716 ( .A(n5424), .Y(n5417) );
  INVX2 U5717 ( .A(n5424), .Y(n5416) );
  INVX2 U5718 ( .A(n1311), .Y(n7178) );
  AND2X1 U5719 ( .A(n7015), .B(n7045), .Y(n2727) );
  INVX2 U5720 ( .A(n2793), .Y(n7319) );
  NAND3X1 U5721 ( .A(n7027), .B(n7034), .C(n7019), .Y(n2601) );
  INVX2 U5722 ( .A(n861), .Y(n7246) );
  NAND2X1 U5723 ( .A(n7328), .B(n7043), .Y(n1826) );
  INVX2 U5724 ( .A(n868), .Y(n7250) );
  INVX2 U5725 ( .A(n211), .Y(n7243) );
  NAND2X1 U5726 ( .A(n2551), .B(n2601), .Y(n2579) );
  INVX2 U5727 ( .A(n2446), .Y(n7309) );
  OR2X1 U5728 ( .A(n5958), .B(n6778), .Y(n6039) );
  INVX2 U5729 ( .A(n5430), .Y(n5458) );
  INVX2 U5730 ( .A(n6992), .Y(n7004) );
  NAND2X1 U5731 ( .A(n7030), .B(n2791), .Y(n2756) );
  NAND4X1 U5732 ( .A(n934), .B(n1993), .C(n6288), .D(n2792), .Y(n2791) );
  AOI222XL U5733 ( .A0(n2710), .A1(n7023), .B0(n7328), .B1(n7319), .C0(n7045), 
        .C1(n7327), .Y(n2792) );
  INVX2 U5734 ( .A(n5430), .Y(n5457) );
  NAND2X1 U5735 ( .A(n5355), .B(n1354), .Y(n1774) );
  INVX2 U5736 ( .A(n1763), .Y(n7218) );
  NOR2X1 U5737 ( .A(n6189), .B(n5384), .Y(n4989) );
  NOR2X1 U5738 ( .A(n6189), .B(n5382), .Y(n4990) );
  INVX2 U5739 ( .A(n6186), .Y(n5384) );
  INVX2 U5740 ( .A(n6090), .Y(n5382) );
  INVX2 U5741 ( .A(n6239), .Y(n7022) );
  NOR2X1 U5742 ( .A(n6189), .B(n5383), .Y(n4991) );
  INVX2 U5743 ( .A(n6719), .Y(n6498) );
  NOR2X1 U5744 ( .A(n2738), .B(n7208), .Y(n2744) );
  NOR2X1 U5745 ( .A(n5389), .B(n6992), .Y(n4992) );
  NAND2BX1 U5746 ( .AN(n2620), .B(n2661), .Y(n2603) );
  NAND2X1 U5747 ( .A(n7197), .B(n1354), .Y(n1859) );
  INVX2 U5748 ( .A(n1848), .Y(n7195) );
  NAND2X1 U5749 ( .A(n7226), .B(n1435), .Y(n1436) );
  NAND2X1 U5750 ( .A(n1354), .B(n4850), .Y(n1457) );
  NAND2X1 U5751 ( .A(n1354), .B(n5351), .Y(n2276) );
  INVX2 U5752 ( .A(n2173), .Y(n7209) );
  BUFX2 U5753 ( .A(n2157), .Y(n5351) );
  OAI31X1 U5754 ( .A0(n7030), .A1(n7034), .A2(n7029), .B0(n7012), .Y(n2157) );
  NOR2X1 U5755 ( .A(n5388), .B(n6992), .Y(n4993) );
  INVX2 U5756 ( .A(n6387), .Y(n5388) );
  NAND2X1 U5757 ( .A(n7219), .B(n1763), .Y(n1746) );
  NAND2X1 U5758 ( .A(n7227), .B(n1381), .Y(n1383) );
  NAND2X1 U5759 ( .A(n1354), .B(n4847), .Y(n1404) );
  INVX2 U5760 ( .A(n2365), .Y(n7203) );
  NOR2X1 U5761 ( .A(n5395), .B(n6992), .Y(n4994) );
  BUFX2 U5762 ( .A(n1995), .Y(n5353) );
  OAI211X1 U5763 ( .A0(n7034), .A1(n7030), .B0(n7019), .C0(n7324), .Y(n1995)
         );
  NAND2X1 U5764 ( .A(n1354), .B(n5353), .Y(n2023) );
  INVX2 U5765 ( .A(n2012), .Y(n7214) );
  NAND2X1 U5766 ( .A(n7210), .B(n2173), .Y(n2156) );
  NOR2X1 U5767 ( .A(n5394), .B(n6992), .Y(n4995) );
  NOR2X1 U5768 ( .A(n5393), .B(n6992), .Y(n4996) );
  NOR2X1 U5769 ( .A(n5392), .B(n6992), .Y(n4997) );
  INVX2 U5770 ( .A(n6716), .Y(n5394) );
  INVX2 U5771 ( .A(n6605), .Y(n5392) );
  INVX2 U5772 ( .A(n6336), .Y(n5387) );
  NAND2X1 U5773 ( .A(n7224), .B(n1536), .Y(n1538) );
  NAND2X1 U5774 ( .A(n1354), .B(n5358), .Y(n1558) );
  NAND2X1 U5775 ( .A(n7222), .B(n1642), .Y(n1643) );
  NAND2X1 U5776 ( .A(n7221), .B(n1691), .Y(n1693) );
  NAND2X1 U5777 ( .A(n1354), .B(n5356), .Y(n1714) );
  NAND2X1 U5778 ( .A(n1354), .B(n5357), .Y(n1662) );
  BUFX2 U5779 ( .A(n1694), .Y(n5356) );
  NAND3X1 U5780 ( .A(n7320), .B(n7030), .C(n7044), .Y(n1694) );
  BUFX2 U5781 ( .A(n1644), .Y(n5357) );
  NAND3X1 U5782 ( .A(n7014), .B(n7030), .C(n7043), .Y(n1644) );
  NAND2X1 U5783 ( .A(n7196), .B(n1848), .Y(n1831) );
  NAND2X1 U5784 ( .A(n7223), .B(n1587), .Y(n1589) );
  NAND2X1 U5785 ( .A(n7225), .B(n1486), .Y(n1488) );
  NAND2X1 U5786 ( .A(n1354), .B(n5359), .Y(n1509) );
  NAND2X1 U5787 ( .A(n1354), .B(n4851), .Y(n1609) );
  NAND2X1 U5788 ( .A(n7213), .B(n1354), .Y(n2102) );
  INVX2 U5789 ( .A(n2091), .Y(n7211) );
  NAND2X1 U5790 ( .A(n7228), .B(n1327), .Y(n1328) );
  NAND2X1 U5791 ( .A(n1354), .B(n5360), .Y(n1351) );
  NOR2X1 U5792 ( .A(n6189), .B(n5385), .Y(n4998) );
  NAND2X1 U5793 ( .A(n7215), .B(n2012), .Y(n1994) );
  INVX2 U5794 ( .A(n6235), .Y(n5385) );
  NAND2X1 U5795 ( .A(n5354), .B(n1354), .Y(n1941) );
  INVX2 U5796 ( .A(n1930), .Y(n7216) );
  INVX2 U5797 ( .A(n739), .Y(n7245) );
  OAI2BB1X1 U5798 ( .A0N(n7015), .A1N(n6498), .B0(n7033), .Y(n6549) );
  NOR2X1 U5799 ( .A(n5391), .B(n6992), .Y(n4999) );
  NOR2X1 U5800 ( .A(n5390), .B(n6992), .Y(n5000) );
  INVX2 U5801 ( .A(n6495), .Y(n5390) );
  INVX2 U5802 ( .A(n2764), .Y(n7205) );
  INVX2 U5803 ( .A(n5949), .Y(n5381) );
  NAND2X1 U5804 ( .A(n7212), .B(n2091), .Y(n2075) );
  NAND2X1 U5805 ( .A(n7217), .B(n1930), .Y(n1913) );
  INVX2 U5806 ( .A(n934), .Y(n7012) );
  AND2X1 U5807 ( .A(n1944), .B(n7034), .Y(n1911) );
  INVX2 U5808 ( .A(n6778), .Y(n6787) );
  NOR2X1 U5809 ( .A(n2743), .B(n7233), .Y(n2750) );
  INVX2 U5810 ( .A(n5402), .Y(n5400) );
  INVX2 U5811 ( .A(n5403), .Y(n5398) );
  INVX2 U5812 ( .A(n5403), .Y(n5399) );
  INVX2 U5813 ( .A(n5402), .Y(n5401) );
  INVX2 U5814 ( .A(n5404), .Y(n5396) );
  INVX2 U5815 ( .A(n5403), .Y(n5397) );
  INVX2 U5816 ( .A(n5433), .Y(n5461) );
  INVX2 U5817 ( .A(n5433), .Y(n5462) );
  INVX2 U5818 ( .A(n5433), .Y(n5463) );
  INVX2 U5819 ( .A(n5428), .Y(n5452) );
  INVX2 U5820 ( .A(n5425), .Y(n5445) );
  INVX2 U5821 ( .A(n5425), .Y(n5443) );
  INVX2 U5822 ( .A(n5429), .Y(n5453) );
  INVX2 U5823 ( .A(n5426), .Y(n5447) );
  INVX2 U5824 ( .A(n5429), .Y(n5454) );
  INVX2 U5825 ( .A(n5427), .Y(n5449) );
  INVX2 U5826 ( .A(n5429), .Y(n5455) );
  INVX2 U5827 ( .A(n5425), .Y(n5444) );
  INVX2 U5828 ( .A(n5430), .Y(n5456) );
  INVX2 U5829 ( .A(n5426), .Y(n5448) );
  INVX2 U5830 ( .A(n5427), .Y(n5450) );
  INVX2 U5831 ( .A(n5427), .Y(n5451) );
  INVX2 U5832 ( .A(n5426), .Y(n5446) );
  INVX2 U5833 ( .A(n5432), .Y(n5460) );
  OAI31XL U5834 ( .A0(n4977), .A1(n5954), .A2(n6028), .B0(n5953), .Y(n5955) );
  AND2X1 U5835 ( .A(n5952), .B(n5951), .Y(n5954) );
  CLKINVXL U5836 ( .A(n6026), .Y(n5953) );
  NOR3BX1 U5837 ( .AN(n2649), .B(n7186), .C(n2650), .Y(n2681) );
  NOR3BX1 U5838 ( .AN(n2681), .B(n2682), .C(n2683), .Y(n2675) );
  NAND3BX1 U5839 ( .AN(n2651), .B(n2647), .C(n2648), .Y(n2650) );
  AND3X2 U5840 ( .A(n7188), .B(n2676), .C(n2675), .Y(n2672) );
  AOI211X1 U5841 ( .A0(n7309), .A1(n7186), .B0(n2620), .C0(n2656), .Y(n2647)
         );
  NOR2X1 U5842 ( .A(n2652), .B(n7177), .Y(n2566) );
  INVX2 U5843 ( .A(n2564), .Y(n7171) );
  NAND2X1 U5844 ( .A(n7186), .B(n7311), .Y(n2648) );
  INVX2 U5845 ( .A(n2563), .Y(n7173) );
  NAND3X1 U5846 ( .A(n2733), .B(n7309), .C(n7187), .Y(n2649) );
  INVX2 U5847 ( .A(n2565), .Y(n7172) );
  AOI2BB1X1 U5848 ( .A0N(n7311), .A1N(n5571), .B0(n7188), .Y(n2682) );
  INVX2 U5849 ( .A(n2680), .Y(n7188) );
  NAND2X1 U5850 ( .A(n2662), .B(n7175), .Y(n2634) );
  AND2X1 U5851 ( .A(n2672), .B(n7187), .Y(n2553) );
  INVX2 U5852 ( .A(n2635), .Y(n7176) );
  AOI222XL U5853 ( .A0(N5132), .A1(n2552), .B0(N5140), .B1(n2553), .C0(N5124), 
        .C1(n2554), .Y(n2616) );
  INVX2 U5854 ( .A(n1585), .Y(n7014) );
  NAND4X1 U5855 ( .A(n2686), .B(n2601), .C(n2661), .D(n2687), .Y(n2656) );
  AOI211X1 U5856 ( .A0(n7030), .A1(n2602), .B0(n2590), .C0(n2591), .Y(n2687)
         );
  INVX2 U5857 ( .A(n2800), .Y(n7328) );
  INVX2 U5858 ( .A(n2805), .Y(n7044) );
  NOR2BX1 U5859 ( .AN(n2675), .B(n2676), .Y(n2554) );
  AND2X1 U5860 ( .A(n2675), .B(n2680), .Y(n2552) );
  AOI222XL U5861 ( .A0(N5118), .A1(n2556), .B0(N5126), .B1(n2554), .C0(N5134), 
        .C1(n2552), .Y(n2587) );
  AOI222XL U5862 ( .A0(n5568), .A1(n2556), .B0(N5125), .B1(n2554), .C0(N5133), 
        .C1(n2552), .Y(n2598) );
  NAND2BX1 U5863 ( .AN(n2106), .B(n7329), .Y(n2723) );
  NOR3X1 U5864 ( .A(n7039), .B(n1743), .C(n7040), .Y(n2710) );
  INVX2 U5865 ( .A(n6552), .Y(n7015) );
  NAND2X1 U5866 ( .A(n7023), .B(n7329), .Y(n2697) );
  INVX2 U5867 ( .A(n2788), .Y(n7023) );
  NAND2X1 U5868 ( .A(n2697), .B(n2704), .Y(n2713) );
  OR2X1 U5869 ( .A(n2106), .B(n7329), .Y(n1864) );
  AND2X1 U5870 ( .A(n2683), .B(n2681), .Y(n2555) );
  AOI222XL U5871 ( .A0(N5094), .A1(n2558), .B0(N5102), .B1(n2557), .C0(N5110), 
        .C1(n2555), .Y(n2586) );
  AOI222XL U5872 ( .A0(N5093), .A1(n2558), .B0(N5101), .B1(n2557), .C0(N5109), 
        .C1(n2555), .Y(n2597) );
  AND2X1 U5873 ( .A(n7186), .B(n2655), .Y(n2568) );
  OAI21X1 U5874 ( .A0(n2446), .A1(n2656), .B0(n2650), .Y(n2655) );
  AOI222XL U5875 ( .A0(N5108), .A1(n2555), .B0(N5061), .B1(n2556), .C0(N5100), 
        .C1(n2557), .Y(n2615) );
  NAND2X1 U5876 ( .A(n7021), .B(n7329), .Y(n2461) );
  INVX2 U5877 ( .A(n1484), .Y(n7016) );
  NOR2X1 U5878 ( .A(n2788), .B(n7329), .Y(n2700) );
  AOI222XL U5879 ( .A0(N5076), .A1(n2567), .B0(N5092), .B1(n2558), .C0(N5068), 
        .C1(n2559), .Y(n2610) );
  AND2X1 U5880 ( .A(n2651), .B(n2647), .Y(n2567) );
  AOI21X1 U5881 ( .A0(n2717), .A1(n7324), .B0(n7031), .Y(n2698) );
  INVX2 U5882 ( .A(n6777), .Y(n7031) );
  NAND2X1 U5883 ( .A(n1827), .B(n7039), .Y(n1863) );
  AOI221XL U5884 ( .A0(n2718), .A1(n1561), .B0(n7043), .B1(n7044), .C0(n7318), 
        .Y(n2638) );
  INVX2 U5885 ( .A(n2720), .Y(n7318) );
  AOI221XL U5886 ( .A0(n2701), .A1(n7013), .B0(n7320), .B1(n2721), .C0(n1944), 
        .Y(n2720) );
  NAND3X1 U5887 ( .A(n5571), .B(n7311), .C(n2680), .Y(n2684) );
  INVX2 U5888 ( .A(n2106), .Y(n7025) );
  NOR2X1 U5889 ( .A(n2800), .B(n2461), .Y(n1944) );
  NAND4X1 U5890 ( .A(n2688), .B(n2630), .C(n2666), .D(n2631), .Y(n2580) );
  NAND2X1 U5891 ( .A(n7031), .B(n7034), .Y(n2688) );
  INVX2 U5892 ( .A(n2689), .Y(n7326) );
  INVX2 U5893 ( .A(n2696), .Y(n7327) );
  INVX2 U5894 ( .A(n2704), .Y(n7320) );
  AND2X1 U5895 ( .A(n2784), .B(n5459), .Y(n2739) );
  OR2X1 U5896 ( .A(n6775), .B(n7329), .Y(n2153) );
  OAI2BB1X1 U5897 ( .A0N(n2689), .A1N(n934), .B0(n7034), .Y(n2631) );
  OR2X1 U5898 ( .A(n2153), .B(n2106), .Y(n934) );
  INVX2 U5899 ( .A(n7230), .Y(n7030) );
  INVX2 U5900 ( .A(n5434), .Y(n5431) );
  AOI2BB1X1 U5901 ( .A0N(n5006), .A1N(n2694), .B0(n6776), .Y(n2668) );
  NOR2X1 U5902 ( .A(n2696), .B(n2697), .Y(n2694) );
  OR2X1 U5903 ( .A(n7028), .B(n2668), .Y(n2590) );
  INVX2 U5904 ( .A(n2735), .Y(n7190) );
  AND2X1 U5905 ( .A(n2784), .B(n5466), .Y(n2737) );
  NAND2X1 U5906 ( .A(n7297), .B(n1290), .Y(n1281) );
  NAND2X1 U5907 ( .A(n7297), .B(n1233), .Y(n1224) );
  NAND3X1 U5908 ( .A(n5571), .B(n1237), .C(n5568), .Y(n1290) );
  NAND2X1 U5909 ( .A(n7297), .B(n1280), .Y(n1271) );
  NAND2X1 U5910 ( .A(n7297), .B(n1247), .Y(n1238) );
  NAND2X1 U5911 ( .A(n7297), .B(n1257), .Y(n1248) );
  OR2X1 U5912 ( .A(n2696), .B(n2723), .Y(n6288) );
  NAND2X1 U5913 ( .A(n7297), .B(n1301), .Y(n1292) );
  NAND2X1 U5914 ( .A(n5568), .B(n1258), .Y(n1301) );
  INVX2 U5915 ( .A(n7206), .Y(n7034) );
  INVX2 U5916 ( .A(n5467), .Y(n5464) );
  NOR2X1 U5917 ( .A(n7035), .B(n2708), .Y(n2716) );
  INVX2 U5918 ( .A(n1233), .Y(n7184) );
  INVX2 U5919 ( .A(n1280), .Y(n7182) );
  INVX2 U5920 ( .A(n1247), .Y(n7183) );
  INVX2 U5921 ( .A(n1257), .Y(n7180) );
  NAND2X1 U5922 ( .A(n7297), .B(n1311), .Y(n1302) );
  NAND2X1 U5923 ( .A(n7297), .B(n1268), .Y(n1259) );
  NAND3X1 U5924 ( .A(n1270), .B(n1269), .C(n5568), .Y(n1311) );
  NAND2X1 U5925 ( .A(n7030), .B(n2724), .Y(n2661) );
  NAND4BX1 U5926 ( .AN(n2072), .B(n1826), .C(n1993), .D(n2725), .Y(n2724) );
  AOI221XL U5927 ( .A0(n7013), .A1(n2721), .B0(n7044), .B1(n7319), .C0(n2727), 
        .Y(n2725) );
  INVX2 U5928 ( .A(n6775), .Y(n7027) );
  OAI2BB2X1 U5929 ( .B0(n7312), .B1(n4848), .A0N(N4595), .A1N(n2376), .Y(n4015) );
  INVX2 U5930 ( .A(n6776), .Y(n7029) );
  INVX2 U5931 ( .A(n117), .Y(n5415) );
  OAI2BB2X1 U5932 ( .B0(n4848), .B1(n7311), .A0N(N4589), .A1N(n2376), .Y(n4021) );
  OAI2BB2X1 U5933 ( .B0(n4848), .B1(n7310), .A0N(N4588), .A1N(n2376), .Y(n4022) );
  INVX2 U5934 ( .A(n7189), .Y(n5423) );
  INVX2 U5935 ( .A(n7189), .Y(n5424) );
  INVX2 U5936 ( .A(n1268), .Y(n7185) );
  OAI2BB2X1 U5937 ( .B0(n7040), .B1(n2354), .A0N(N4699), .A1N(n7042), .Y(n3995) );
  OAI2BB2X1 U5938 ( .B0(n7329), .B1(n2354), .A0N(N4697), .A1N(n7042), .Y(n3997) );
  OAI2BB2X1 U5939 ( .B0(n7039), .B1(n2354), .A0N(N4696), .A1N(n7042), .Y(n3998) );
  OAI211X1 U5940 ( .A0(n761), .A1(n7427), .B0(n774), .C0(n775), .Y(n186) );
  NAND2X1 U5941 ( .A(N9759), .B(n7275), .Y(n774) );
  INVX2 U5942 ( .A(N9710), .Y(n7427) );
  AOI222XL U5943 ( .A0(N9857), .A1(n7286), .B0(N9906), .B1(n7264), .C0(N9808), 
        .C1(n7277), .Y(n775) );
  NOR2X1 U5944 ( .A(n1779), .B(n2700), .Y(n2793) );
  AOI21X1 U5945 ( .A0(n2728), .A1(n2729), .B0(n7230), .Y(n2620) );
  AOI211X1 U5946 ( .A0(n7015), .A1(n7013), .B0(n2730), .C0(n2731), .Y(n2729)
         );
  AOI222XL U5947 ( .A0(n1561), .A1(n7046), .B0(n7016), .B1(n7032), .C0(n2710), 
        .C1(n7319), .Y(n2728) );
  NOR2X1 U5948 ( .A(n5363), .B(n272), .Y(n346) );
  AND4X2 U5949 ( .A(n822), .B(n407), .C(n851), .D(n852), .Y(n198) );
  NOR3X1 U5950 ( .A(n719), .B(n718), .C(n720), .Y(n851) );
  NOR4X1 U5951 ( .A(n777), .B(n821), .C(n815), .D(n814), .Y(n852) );
  NAND4BBX1 U5952 ( .AN(n591), .BN(n589), .C(n871), .D(n872), .Y(n821) );
  AOI21X1 U5953 ( .A0(n7279), .A1(n869), .B0(n714), .Y(n871) );
  AOI211X1 U5954 ( .A0(n5015), .A1(n870), .B0(n590), .C0(n715), .Y(n872) );
  BUFX2 U5955 ( .A(n180), .Y(n5363) );
  NAND4X1 U5956 ( .A(n198), .B(n816), .C(n343), .D(n802), .Y(n180) );
  NOR3BX1 U5957 ( .AN(n877), .B(n765), .C(n764), .Y(n739) );
  NOR2X1 U5958 ( .A(n869), .B(n7255), .Y(n861) );
  AOI2BB2X1 U5959 ( .B0(n7246), .B1(n7261), .A0N(n921), .A1N(n802), .Y(n877)
         );
  NOR2X1 U5960 ( .A(n7246), .B(n857), .Y(n921) );
  OR2X1 U5961 ( .A(n918), .B(n7257), .Y(n869) );
  NOR2X1 U5962 ( .A(n5363), .B(n831), .Y(n279) );
  INVX2 U5963 ( .A(n928), .Y(n7258) );
  NOR2X1 U5964 ( .A(n1585), .B(n2723), .Y(n2731) );
  NAND2X1 U5965 ( .A(n853), .B(n854), .Y(n814) );
  AOI222XL U5966 ( .A0(n7257), .A1(n7281), .B0(n7272), .B1(n857), .C0(n7260), 
        .C1(n7281), .Y(n853) );
  AOI221XL U5967 ( .A0(n7272), .A1(n7246), .B0(n7265), .B1(n857), .C0(n721), 
        .Y(n854) );
  OR2X1 U5968 ( .A(n186), .B(n197), .Y(n742) );
  INVX2 U5969 ( .A(n295), .Y(n6956) );
  NOR2BX1 U5970 ( .AN(n199), .B(n5363), .Y(n464) );
  NOR2X1 U5971 ( .A(n867), .B(n861), .Y(n812) );
  NOR2X1 U5972 ( .A(n1484), .B(n2788), .Y(n2730) );
  NOR2X1 U5973 ( .A(n5363), .B(n182), .Y(n211) );
  NOR2X1 U5974 ( .A(n5363), .B(n169), .Y(n600) );
  INVX2 U5975 ( .A(n884), .Y(n7264) );
  AOI222XL U5976 ( .A0(n857), .A1(n7275), .B0(n918), .B1(n7286), .C0(n7244), 
        .C1(n7264), .Y(n862) );
  INVX2 U5977 ( .A(n178), .Y(n7281) );
  INVX2 U5978 ( .A(n182), .Y(n7265) );
  INVX2 U5979 ( .A(n272), .Y(n7279) );
  INVX2 U5980 ( .A(n882), .Y(n7286) );
  NAND2X1 U5981 ( .A(n7265), .B(n7244), .Y(n584) );
  INVX2 U5982 ( .A(n301), .Y(n6958) );
  INVX2 U5983 ( .A(n761), .Y(n7261) );
  NOR2X1 U5984 ( .A(n5363), .B(n178), .Y(n598) );
  NOR2X1 U5985 ( .A(n870), .B(n7257), .Y(n868) );
  INVX2 U5986 ( .A(n857), .Y(n7251) );
  INVX2 U5987 ( .A(n359), .Y(n6932) );
  INVX2 U5988 ( .A(n416), .Y(n6908) );
  NAND2X1 U5989 ( .A(n7249), .B(n199), .Y(n586) );
  INVX2 U5990 ( .A(n2494), .Y(n7291) );
  INVX2 U5991 ( .A(n422), .Y(n6910) );
  INVX2 U5992 ( .A(n365), .Y(n6934) );
  AOI22X1 U5993 ( .A0(n7260), .A1(n7264), .B0(n7250), .B1(n7286), .Y(n823) );
  AOI21X1 U5994 ( .A0(N9710), .A1(n7261), .B0(n197), .Y(n737) );
  INVX2 U5995 ( .A(n867), .Y(n7277) );
  AND4X2 U5996 ( .A(n182), .B(n831), .C(n838), .D(n839), .Y(n185) );
  NOR3X1 U5997 ( .A(n7290), .B(n5015), .C(n7281), .Y(n838) );
  NOR4X1 U5998 ( .A(n7272), .B(n199), .C(n7279), .D(n840), .Y(n839) );
  INVX2 U5999 ( .A(n610), .Y(n6836) );
  NOR4BBX1 U6000 ( .AN(n592), .BN(n594), .C(n344), .D(n597), .Y(n816) );
  INVX2 U6001 ( .A(n831), .Y(n7267) );
  NAND2X1 U6002 ( .A(n7267), .B(n7257), .Y(n594) );
  AOI21X1 U6003 ( .A0(n2602), .A1(n7030), .B0(n2603), .Y(n2551) );
  NAND2X1 U6004 ( .A(n7267), .B(n7255), .Y(n592) );
  NAND2X1 U6005 ( .A(n7290), .B(n7254), .Y(n407) );
  INVX2 U6006 ( .A(n169), .Y(n7290) );
  AOI22X1 U6007 ( .A0(n869), .A1(n7290), .B0(n870), .B1(n7281), .Y(n822) );
  INVX2 U6008 ( .A(n476), .Y(n6884) );
  INVX2 U6009 ( .A(n532), .Y(n6860) );
  INVX2 U6010 ( .A(n616), .Y(n6838) );
  INVX2 U6011 ( .A(n225), .Y(n6975) );
  INVX2 U6012 ( .A(n224), .Y(n6977) );
  NAND2X1 U6013 ( .A(n7267), .B(n7249), .Y(n343) );
  INVX2 U6014 ( .A(n666), .Y(n6812) );
  INVX2 U6015 ( .A(n229), .Y(n6979) );
  INVX2 U6016 ( .A(n227), .Y(n6980) );
  INVX2 U6017 ( .A(n734), .Y(n7041) );
  INVX2 U6018 ( .A(n672), .Y(n6814) );
  INVX2 U6019 ( .A(n668), .Y(n6803) );
  INVX2 U6020 ( .A(n671), .Y(n6816) );
  INVX2 U6021 ( .A(n538), .Y(n6862) );
  INVX2 U6022 ( .A(n482), .Y(n6886) );
  NAND2X1 U6023 ( .A(n7310), .B(n7311), .Y(n2446) );
  OAI31X1 U6024 ( .A0(n2794), .A1(n7328), .A2(n1907), .B0(n7030), .Y(n2757) );
  NAND3BX1 U6025 ( .AN(n5013), .B(n2696), .C(n7323), .Y(n2794) );
  NAND4BBX1 U6026 ( .AN(n814), .BN(n815), .C(n816), .D(n817), .Y(n785) );
  NOR3X1 U6027 ( .A(n818), .B(n819), .C(n7247), .Y(n817) );
  OR2X1 U6028 ( .A(n5458), .B(n5465), .Y(n5895) );
  OR2X1 U6029 ( .A(n5001), .B(n6030), .Y(n6778) );
  NOR2X1 U6030 ( .A(n5412), .B(n6790), .Y(n5001) );
  INVX2 U6031 ( .A(n5001), .Y(n1354) );
  INVX2 U6032 ( .A(n6037), .Y(n5958) );
  INVX2 U6033 ( .A(n7007), .Y(n5412) );
  INVX2 U6034 ( .A(n5435), .Y(n5430) );
  OR2X1 U6035 ( .A(n5350), .B(n5442), .Y(n6992) );
  NAND4X1 U6036 ( .A(n2762), .B(n2763), .C(n2796), .D(n2774), .Y(n2754) );
  OAI2BB1X1 U6037 ( .A0N(n2801), .A1N(n2802), .B0(n7030), .Y(n2763) );
  AOI221XL U6038 ( .A0(n2710), .A1(n7013), .B0(n7043), .B1(n7015), .C0(n2730), 
        .Y(n2802) );
  AOI222XL U6039 ( .A0(n7324), .A1(n1561), .B0(n7044), .B1(n7021), .C0(n7320), 
        .C1(n7046), .Y(n2801) );
  OAI211X1 U6040 ( .A0(n2776), .A1(n7230), .B0(n2807), .C0(n2766), .Y(n2795)
         );
  INVX2 U6041 ( .A(n917), .Y(n7247) );
  AOI211X1 U6042 ( .A0(n918), .A1(n7275), .B0(n765), .C0(n764), .Y(n917) );
  NAND3X1 U6043 ( .A(n5352), .B(n7264), .C(n7219), .Y(n1763) );
  BUFX2 U6044 ( .A(n1747), .Y(n5355) );
  AOI33X1 U6045 ( .A0(n7328), .A1(n7034), .A2(n1779), .B0(n1779), .B1(n7030), 
        .B2(n7044), .Y(n1747) );
  NOR2X1 U6046 ( .A(n5350), .B(n5386), .Y(n5002) );
  OAI221X1 U6047 ( .A0(n6792), .A1(n1863), .B0(n1988), .B1(n7206), .C0(n6140), 
        .Y(n6186) );
  AOI221XL U6048 ( .A0(n7326), .A1(n7023), .B0(n7324), .B1(n7019), .C0(n7317), 
        .Y(n1988) );
  AOI31X1 U6049 ( .A0(n1827), .A1(n7030), .A2(n7045), .B0(n5350), .Y(n6140) );
  OAI221X1 U6050 ( .A0(n6044), .A1(n6719), .B0(n1826), .B1(n7206), .C0(n6043), 
        .Y(n6090) );
  AOI2BB1X1 U6051 ( .A0N(n2106), .A1N(n6042), .B0(n7328), .Y(n6044) );
  AOI31X1 U6052 ( .A0(n1829), .A1(n7030), .A2(n7044), .B0(n5350), .Y(n6043) );
  INVX2 U6053 ( .A(n1827), .Y(n6042) );
  INVX2 U6054 ( .A(n6286), .Y(n5386) );
  OR2X1 U6055 ( .A(n2153), .B(n2788), .Y(n6239) );
  OR2X1 U6056 ( .A(n7230), .B(n7329), .Y(n6719) );
  INVX2 U6057 ( .A(n6138), .Y(n5383) );
  NAND4BX1 U6058 ( .AN(n2754), .B(n2755), .C(n2756), .D(n2757), .Y(n2738) );
  NAND2X1 U6059 ( .A(n7030), .B(n2758), .Y(n2755) );
  OR2X1 U6060 ( .A(n1484), .B(n7230), .Y(n6444) );
  INVX2 U6061 ( .A(n6441), .Y(n5389) );
  INVX2 U6062 ( .A(n1862), .Y(n7197) );
  OAI32X1 U6063 ( .A0(n1863), .A1(n1864), .A2(n7230), .B0(n7206), .B1(n1826), 
        .Y(n1862) );
  NAND3X1 U6064 ( .A(n5352), .B(n7286), .C(n7196), .Y(n1848) );
  NAND3X1 U6065 ( .A(n5352), .B(n7281), .C(n7226), .Y(n1435) );
  NAND3X1 U6066 ( .A(n5352), .B(n7285), .C(n7210), .Y(n2173) );
  NAND2BX1 U6067 ( .AN(n5350), .B(n4847), .Y(n6387) );
  OR2X1 U6068 ( .A(n7230), .B(n6793), .Y(n6391) );
  INVX2 U6069 ( .A(n889), .Y(n7003) );
  AOI211X1 U6070 ( .A0(n890), .A1(n743), .B0(n7282), .C0(n812), .Y(n889) );
  OR2X1 U6071 ( .A(n835), .B(n7047), .Y(n890) );
  NAND3X1 U6072 ( .A(n5352), .B(n7290), .C(n7227), .Y(n1381) );
  INVX2 U6073 ( .A(n5350), .Y(n7033) );
  NAND2X1 U6074 ( .A(n7033), .B(n7297), .Y(n2365) );
  INVX2 U6075 ( .A(n6771), .Y(n5395) );
  INVX2 U6076 ( .A(n777), .Y(n6984) );
  NAND3X1 U6077 ( .A(n5352), .B(n7275), .C(n7215), .Y(n2012) );
  OAI211X1 U6078 ( .A0(n6721), .A1(n6719), .B0(n6665), .C0(n7033), .Y(n6716)
         );
  OAI211X1 U6079 ( .A0(n1585), .A1(n6719), .B0(n4851), .C0(n7033), .Y(n6605)
         );
  INVX2 U6080 ( .A(n6661), .Y(n5393) );
  INVX2 U6081 ( .A(n6774), .Y(n7020) );
  NAND4BX1 U6082 ( .AN(n719), .B(n407), .C(n343), .D(n811), .Y(n786) );
  NOR4X1 U6083 ( .A(n812), .B(n7282), .C(n718), .D(n720), .Y(n811) );
  NOR2X1 U6084 ( .A(n5350), .B(n5387), .Y(n5003) );
  NAND3X1 U6085 ( .A(n6290), .B(n7033), .C(n6289), .Y(n6336) );
  OAI2BB1X1 U6086 ( .A0N(n6774), .A1N(n6288), .B0(n7034), .Y(n6290) );
  OAI2BB1X1 U6087 ( .A0N(n7230), .A1N(n6776), .B0(n6987), .Y(n6289) );
  NAND3X1 U6088 ( .A(n5352), .B(n7265), .C(n7224), .Y(n1536) );
  BUFX2 U6089 ( .A(n1539), .Y(n5358) );
  NAND3X1 U6090 ( .A(n7015), .B(n7030), .C(n1561), .Y(n1539) );
  NAND3X1 U6091 ( .A(n5352), .B(n5015), .C(n7221), .Y(n1691) );
  NAND3X1 U6092 ( .A(n5352), .B(n7279), .C(n7222), .Y(n1642) );
  NOR2X1 U6093 ( .A(n840), .B(n7285), .Y(n743) );
  NAND3X1 U6094 ( .A(n5352), .B(n199), .C(n7223), .Y(n1587) );
  NAND3X1 U6095 ( .A(n5352), .B(n7272), .C(n7225), .Y(n1486) );
  INVX2 U6096 ( .A(n2105), .Y(n7213) );
  OAI22X1 U6097 ( .A0(n2106), .A1(n2070), .B0(n2107), .B1(n2108), .Y(n2105) );
  NOR2X1 U6098 ( .A(n7034), .B(n7029), .Y(n2107) );
  NAND3X1 U6099 ( .A(n5352), .B(n7261), .C(n7212), .Y(n2091) );
  NAND2BX1 U6100 ( .AN(n7230), .B(n7326), .Y(n2070) );
  BUFX2 U6101 ( .A(n1489), .Y(n5359) );
  NAND3X1 U6102 ( .A(n7030), .B(n7021), .C(n7016), .Y(n1489) );
  NAND3X1 U6103 ( .A(n7228), .B(n7267), .C(n5352), .Y(n1327) );
  BUFX2 U6104 ( .A(n1329), .Y(n5360) );
  NAND3X1 U6105 ( .A(n7030), .B(n7032), .C(n7017), .Y(n1329) );
  INVX2 U6106 ( .A(n6793), .Y(n7017) );
  INVX2 U6107 ( .A(n802), .Y(n7285) );
  NAND3BX1 U6108 ( .AN(n5350), .B(n2070), .C(n5004), .Y(n6235) );
  NAND2X1 U6109 ( .A(n6188), .B(n7034), .Y(n5004) );
  NAND3X1 U6110 ( .A(n5352), .B(n7277), .C(n7217), .Y(n1930) );
  INVX2 U6111 ( .A(n6041), .Y(n6189) );
  OAI2BB1X1 U6112 ( .A0N(n5466), .A1N(n7033), .B0(n6992), .Y(n6041) );
  OAI2BB1X1 U6113 ( .A0N(n6445), .A1N(n2106), .B0(n7033), .Y(n6495) );
  INVX2 U6114 ( .A(n6444), .Y(n6445) );
  NAND2X1 U6115 ( .A(n2772), .B(n7032), .Y(n2764) );
  NOR2X1 U6116 ( .A(n5350), .B(n5381), .Y(n5005) );
  OR2X1 U6117 ( .A(n5350), .B(n6030), .Y(n5949) );
  INVX2 U6118 ( .A(n1350), .Y(n7269) );
  NAND2X1 U6119 ( .A(n7034), .B(n2808), .Y(n2766) );
  OAI2BB1X1 U6120 ( .A0N(n2701), .A1N(n7013), .B0(n2696), .Y(n2808) );
  OR2X1 U6121 ( .A(n5350), .B(n6993), .Y(n7002) );
  OR2X1 U6122 ( .A(n7018), .B(n5013), .Y(n6987) );
  BUFX2 U6123 ( .A(n1914), .Y(n5354) );
  AOI2BB1X1 U6124 ( .A0N(n1826), .A1N(n7230), .B0(n1911), .Y(n1914) );
  INVX2 U6125 ( .A(n2265), .Y(n5901) );
  AND2X1 U6126 ( .A(n1779), .B(n7324), .Y(n2073) );
  INVX2 U6127 ( .A(n2022), .Y(n7274) );
  INVX2 U6128 ( .A(n7121), .Y(n7124) );
  INVX2 U6129 ( .A(n1661), .Y(n7278) );
  INVX2 U6130 ( .A(n1940), .Y(n7276) );
  NAND3X1 U6131 ( .A(n2764), .B(n2765), .C(n2766), .Y(n2743) );
  INVX2 U6132 ( .A(n1608), .Y(n7288) );
  AND2X1 U6133 ( .A(n2796), .B(n2807), .Y(n2768) );
  INVX2 U6134 ( .A(n1508), .Y(n7271) );
  NAND3X1 U6135 ( .A(n2763), .B(n2774), .C(n2764), .Y(n2773) );
  INVX2 U6136 ( .A(n6030), .Y(n6035) );
  INVX2 U6137 ( .A(n7007), .Y(n5413) );
  INVX2 U6138 ( .A(n7007), .Y(n5411) );
  INVX2 U6139 ( .A(n7007), .Y(n5410) );
  INVX2 U6140 ( .A(n7007), .Y(n5409) );
  INVX2 U6141 ( .A(n7007), .Y(n5408) );
  INVX2 U6142 ( .A(n7007), .Y(n5407) );
  INVX2 U6143 ( .A(n7007), .Y(n5406) );
  INVX2 U6144 ( .A(n7007), .Y(n5405) );
  INVX2 U6145 ( .A(n7007), .Y(n5402) );
  INVX2 U6146 ( .A(n7007), .Y(n5414) );
  INVX2 U6147 ( .A(n7007), .Y(n5403) );
  OAI2BB1X1 U6148 ( .A0N(n7021), .A1N(n2772), .B0(n2756), .Y(n2781) );
  INVX2 U6149 ( .A(n6664), .Y(n6721) );
  OAI31X1 U6150 ( .A0(n1743), .A1(n7040), .A2(n7035), .B0(n7323), .Y(n6664) );
  INVX2 U6151 ( .A(n7007), .Y(n5404) );
  AOI33X1 U6152 ( .A0(n2436), .A1(n7308), .A2(n2445), .B0(n2454), .B1(n2446), 
        .B2(N5059), .Y(n2453) );
  AOI221XL U6153 ( .A0(n2449), .A1(n7306), .B0(n2451), .B1(n2433), .C0(n7220), 
        .Y(WEN13) );
  INVX2 U6154 ( .A(n2456), .Y(n7306) );
  NOR2X1 U6155 ( .A(n2432), .B(n2442), .Y(n2451) );
  INVX2 U6156 ( .A(n2453), .Y(n7220) );
  AOI222XL U6157 ( .A0(n2435), .A1(n7300), .B0(n2456), .B1(n2449), .C0(n2454), 
        .C1(n2448), .Y(WEN03) );
  INVX2 U6158 ( .A(n2430), .Y(n7308) );
  OAI211X1 U6159 ( .A0(n5568), .A1(n7307), .B0(n2428), .C0(n2429), .Y(WEN73)
         );
  OAI2BB1X1 U6160 ( .A0N(n2430), .A1N(n1270), .B0(n5568), .Y(n2428) );
  AND2X1 U6161 ( .A(n2433), .B(n7301), .Y(n2429) );
  NAND4X1 U6162 ( .A(n2431), .B(n2429), .C(n5568), .D(N5061), .Y(WEN63) );
  NAND3BX1 U6163 ( .AN(n2432), .B(n5568), .C(n2429), .Y(WEN53) );
  NAND3X1 U6164 ( .A(n5568), .B(n7301), .C(n2435), .Y(WEN43) );
  INVX2 U6165 ( .A(n2439), .Y(n7301) );
  OAI211X1 U6166 ( .A0(n835), .A1(n7047), .B0(n761), .C0(n802), .Y(n874) );
  INVX2 U6167 ( .A(n1456), .Y(n7280) );
  INVX2 U6168 ( .A(n2272), .Y(n7284) );
  XOR2X1 U6169 ( .A(n2430), .B(n5571), .Y(n2431) );
  INVX2 U6170 ( .A(n1455), .Y(n7507) );
  INVX2 U6171 ( .A(n5434), .Y(n5433) );
  NAND2X1 U6172 ( .A(N5061), .B(n5571), .Y(n2440) );
  INVX2 U6173 ( .A(n104), .Y(n7307) );
  INVX2 U6174 ( .A(n2442), .Y(n7300) );
  AOI2BB1X1 U6175 ( .A0N(n7310), .A1N(n7311), .B0(n7309), .Y(n2456) );
  OR2X1 U6176 ( .A(n5458), .B(n5465), .Y(n5349) );
  OR2X1 U6177 ( .A(n5458), .B(n5465), .Y(n5348) );
  INVX2 U6178 ( .A(n5435), .Y(n5428) );
  INVX2 U6179 ( .A(n5435), .Y(n5429) );
  INVX2 U6180 ( .A(n5436), .Y(n5425) );
  INVX2 U6181 ( .A(n5436), .Y(n5427) );
  INVX2 U6182 ( .A(n5436), .Y(n5426) );
  INVX2 U6183 ( .A(n5434), .Y(n5432) );
  OR2X1 U6184 ( .A(n6913), .B(n6716), .Y(n6667) );
  OR2X1 U6185 ( .A(n6966), .B(n6605), .Y(n6555) );
  OR2X1 U6186 ( .A(n6865), .B(n6661), .Y(n6611) );
  OR2X1 U6187 ( .A(n6889), .B(n6771), .Y(n6723) );
  OAI2BB1X1 U6188 ( .A0N(N6291), .A1N(n4996), .B0(n6610), .Y(n3467) );
  OR2X1 U6189 ( .A(n6859), .B(n6661), .Y(n6610) );
  OR2X1 U6190 ( .A(n6817), .B(n6495), .Y(n6447) );
  OR2X1 U6191 ( .A(n6841), .B(n6441), .Y(n6393) );
  OR2X1 U6192 ( .A(n6937), .B(n6549), .Y(n6500) );
  OR2X1 U6193 ( .A(n6954), .B(n6387), .Y(n6339) );
  OR2X1 U6194 ( .A(n6907), .B(n6716), .Y(n6666) );
  OR2X1 U6195 ( .A(n6883), .B(n6771), .Y(n6722) );
  OR2X1 U6196 ( .A(n6911), .B(n6716), .Y(n6668) );
  OR2X1 U6197 ( .A(n6965), .B(n6605), .Y(n6556) );
  OR2X1 U6198 ( .A(n6835), .B(n6441), .Y(n6392) );
  OR2X1 U6199 ( .A(n6951), .B(n6387), .Y(n6338) );
  OR2X1 U6200 ( .A(n6931), .B(n6549), .Y(n6499) );
  OR2X1 U6201 ( .A(n6863), .B(n6661), .Y(n6612) );
  OAI2BB1X1 U6202 ( .A0N(N6285), .A1N(n4996), .B0(n6617), .Y(n3473) );
  OR2X1 U6203 ( .A(n6857), .B(n6661), .Y(n6617) );
  OR2X1 U6204 ( .A(n6858), .B(n6661), .Y(n6616) );
  OR2X1 U6205 ( .A(n6811), .B(n6495), .Y(n6446) );
  OR2X1 U6206 ( .A(n6968), .B(n6605), .Y(n6568) );
  OAI2BB1X1 U6207 ( .A0N(N6244), .A1N(n4995), .B0(n6673), .Y(n3528) );
  OR2X1 U6208 ( .A(n6905), .B(n6716), .Y(n6673) );
  OR2X1 U6209 ( .A(n6906), .B(n6716), .Y(n6672) );
  OR2X1 U6210 ( .A(n6866), .B(n6771), .Y(n6735) );
  OR2X1 U6211 ( .A(n6915), .B(n6549), .Y(n6511) );
  OAI2BB1X1 U6212 ( .A0N(N6367), .A1N(n4999), .B0(n6506), .Y(n3363) );
  OR2X1 U6213 ( .A(n6929), .B(n6549), .Y(n6506) );
  OR2X1 U6214 ( .A(n6930), .B(n6549), .Y(n6505) );
  OR2X1 U6215 ( .A(n6935), .B(n6549), .Y(n6501) );
  OAI2BB1X1 U6216 ( .A0N(N6326), .A1N(n4997), .B0(n6562), .Y(n3418) );
  OR2X1 U6217 ( .A(n6962), .B(n6605), .Y(n6562) );
  OR2X1 U6218 ( .A(n6963), .B(n6605), .Y(n6561) );
  OR2X1 U6219 ( .A(n6815), .B(n6495), .Y(n6448) );
  OR2X1 U6220 ( .A(n6839), .B(n6441), .Y(n6394) );
  OR2X1 U6221 ( .A(n6953), .B(n6387), .Y(n6340) );
  OR2X1 U6222 ( .A(n6833), .B(n6441), .Y(n6399) );
  OR2X1 U6223 ( .A(n6834), .B(n6441), .Y(n6398) );
  OR2X1 U6224 ( .A(n6959), .B(n6387), .Y(n6345) );
  OR2X1 U6225 ( .A(n6961), .B(n6387), .Y(n6344) );
  OR2X1 U6226 ( .A(n6914), .B(n6549), .Y(n6512) );
  OR2X1 U6227 ( .A(n6809), .B(n6495), .Y(n6453) );
  OR2X1 U6228 ( .A(n6810), .B(n6495), .Y(n6452) );
  OR2X1 U6229 ( .A(n6887), .B(n6771), .Y(n6724) );
  OR2X1 U6230 ( .A(n6855), .B(n6661), .Y(n6615) );
  OR2X1 U6231 ( .A(n6903), .B(n6716), .Y(n6671) );
  OR2X1 U6232 ( .A(n6867), .B(n6771), .Y(n6734) );
  OR2X1 U6233 ( .A(n6882), .B(n6771), .Y(n6728) );
  OAI2BB1X1 U6234 ( .A0N(N6369), .A1N(n4999), .B0(n6504), .Y(n3361) );
  OR2X1 U6235 ( .A(n6927), .B(n6549), .Y(n6504) );
  OR2X1 U6236 ( .A(n6831), .B(n6441), .Y(n6397) );
  OR2X1 U6237 ( .A(n6955), .B(n6387), .Y(n6343) );
  OAI2BB1X1 U6238 ( .A0N(N6203), .A1N(n4994), .B0(n6729), .Y(n3583) );
  OR2X1 U6239 ( .A(n6881), .B(n6771), .Y(n6729) );
  OR2X1 U6240 ( .A(n6807), .B(n6495), .Y(n6451) );
  OR2X1 U6241 ( .A(n6939), .B(n6387), .Y(n6350) );
  OR2X1 U6242 ( .A(n6938), .B(n6387), .Y(n6351) );
  OR2X1 U6243 ( .A(n6969), .B(n6605), .Y(n6567) );
  OR2X1 U6244 ( .A(n6891), .B(n6716), .Y(n6678) );
  OR2X1 U6245 ( .A(n6890), .B(n6716), .Y(n6679) );
  OR2X1 U6246 ( .A(n6879), .B(n6771), .Y(n6727) );
  OR2X1 U6247 ( .A(n6818), .B(n6441), .Y(n6405) );
  OR2X1 U6248 ( .A(n6794), .B(n6495), .Y(n6459) );
  OR2X1 U6249 ( .A(n6842), .B(n6661), .Y(n6623) );
  OR2X1 U6250 ( .A(n6819), .B(n6441), .Y(n6404) );
  OR2X1 U6251 ( .A(n6843), .B(n6661), .Y(n6622) );
  OR2X1 U6252 ( .A(n6795), .B(n6495), .Y(n6458) );
  OR2X1 U6253 ( .A(n6894), .B(n6716), .Y(n6684) );
  OAI2BB1X1 U6254 ( .A0N(N6236), .A1N(n4995), .B0(n6685), .Y(n3536) );
  OR2X1 U6255 ( .A(n6893), .B(n6716), .Y(n6685) );
  OAI2BB1X1 U6256 ( .A0N(N6441), .A1N(n4992), .B0(n6411), .Y(n3261) );
  OR2X1 U6257 ( .A(n6821), .B(n6441), .Y(n6411) );
  OR2X1 U6258 ( .A(n6822), .B(n6441), .Y(n6410) );
  OAI2BB1X1 U6259 ( .A0N(N6277), .A1N(n4996), .B0(n6629), .Y(n3481) );
  OR2X1 U6260 ( .A(n6845), .B(n6661), .Y(n6629) );
  OR2X1 U6261 ( .A(n6846), .B(n6661), .Y(n6628) );
  OR2X1 U6262 ( .A(n6972), .B(n6605), .Y(n6572) );
  OAI2BB1X1 U6263 ( .A0N(N6400), .A1N(n5000), .B0(n6465), .Y(n3316) );
  OR2X1 U6264 ( .A(n6797), .B(n6495), .Y(n6465) );
  OR2X1 U6265 ( .A(n6798), .B(n6495), .Y(n6464) );
  OAI2BB1X1 U6266 ( .A0N(N6318), .A1N(n4997), .B0(n6573), .Y(n3426) );
  OR2X1 U6267 ( .A(n6971), .B(n6605), .Y(n6573) );
  OR2X1 U6268 ( .A(n6870), .B(n6771), .Y(n6739) );
  OR2X1 U6269 ( .A(n6917), .B(n6549), .Y(n6517) );
  OAI2BB1X1 U6270 ( .A0N(N6360), .A1N(n4999), .B0(n6516), .Y(n3370) );
  OR2X1 U6271 ( .A(n6918), .B(n6549), .Y(n6516) );
  OAI2BB1X1 U6272 ( .A0N(N6195), .A1N(n4994), .B0(n6740), .Y(n3591) );
  OR2X1 U6273 ( .A(n6869), .B(n6771), .Y(n6740) );
  OAI2BB1X1 U6274 ( .A0N(N6482), .A1N(n4993), .B0(n6357), .Y(n3206) );
  OR2X1 U6275 ( .A(n6941), .B(n6387), .Y(n6357) );
  OR2X1 U6276 ( .A(n6942), .B(n6387), .Y(n6356) );
  OAI2BB1X1 U6277 ( .A0N(N6192), .A1N(n4994), .B0(n6744), .Y(n3594) );
  OR2X1 U6278 ( .A(n6873), .B(n6771), .Y(n6744) );
  OR2X1 U6279 ( .A(n6897), .B(n6716), .Y(n6689) );
  OR2X1 U6280 ( .A(n6896), .B(n6716), .Y(n6690) );
  OAI2BB1X1 U6281 ( .A0N(N6315), .A1N(n4997), .B0(n6578), .Y(n3429) );
  OR2X1 U6282 ( .A(n6976), .B(n6605), .Y(n6578) );
  OR2X1 U6283 ( .A(n6849), .B(n6661), .Y(n6634) );
  OAI2BB1X1 U6284 ( .A0N(N6356), .A1N(n4999), .B0(n6522), .Y(n3374) );
  OR2X1 U6285 ( .A(n6921), .B(n6549), .Y(n6522) );
  OAI2BB1X1 U6286 ( .A0N(N6396), .A1N(n5000), .B0(n6469), .Y(n3320) );
  OR2X1 U6287 ( .A(n6800), .B(n6495), .Y(n6469) );
  OAI2BB1X1 U6288 ( .A0N(N6191), .A1N(n4994), .B0(n6745), .Y(n3595) );
  OR2X1 U6289 ( .A(n6872), .B(n6771), .Y(n6745) );
  OAI2BB1X1 U6290 ( .A0N(N6397), .A1N(n5000), .B0(n6468), .Y(n3319) );
  OR2X1 U6291 ( .A(n6801), .B(n6495), .Y(n6468) );
  OAI2BB1X1 U6292 ( .A0N(N6438), .A1N(n4992), .B0(n6414), .Y(n3264) );
  OR2X1 U6293 ( .A(n6825), .B(n6441), .Y(n6414) );
  OAI2BB1X1 U6294 ( .A0N(N6479), .A1N(n4993), .B0(n6360), .Y(n3209) );
  OR2X1 U6295 ( .A(n6945), .B(n6387), .Y(n6360) );
  OAI2BB1X1 U6296 ( .A0N(N6314), .A1N(n4997), .B0(n6579), .Y(n3430) );
  OR2X1 U6297 ( .A(n6974), .B(n6605), .Y(n6579) );
  OAI2BB1X1 U6298 ( .A0N(N6231), .A1N(n4995), .B0(n6691), .Y(n3541) );
  OR2X1 U6299 ( .A(n4865), .B(n6716), .Y(n6691) );
  OR2X1 U6300 ( .A(n6920), .B(n6549), .Y(n6523) );
  OAI2BB1X1 U6301 ( .A0N(N6273), .A1N(n4996), .B0(n6635), .Y(n3485) );
  OR2X1 U6302 ( .A(n6848), .B(n6661), .Y(n6635) );
  OAI2BB1X1 U6303 ( .A0N(N6436), .A1N(n4992), .B0(n6416), .Y(n3266) );
  OR2X1 U6304 ( .A(n4884), .B(n6441), .Y(n6416) );
  OAI2BB1X1 U6305 ( .A0N(N6437), .A1N(n4992), .B0(n6415), .Y(n3265) );
  OR2X1 U6306 ( .A(n6824), .B(n6441), .Y(n6415) );
  OAI2BB1X1 U6307 ( .A0N(N6354), .A1N(n4999), .B0(n6524), .Y(n3376) );
  OR2X1 U6308 ( .A(n4854), .B(n6549), .Y(n6524) );
  OAI2BB1X1 U6309 ( .A0N(N6230), .A1N(n4995), .B0(n6692), .Y(n3542) );
  OR2X1 U6310 ( .A(n4916), .B(n6716), .Y(n6692) );
  NOR3BX1 U6311 ( .AN(N5018), .B(n2652), .C(n1313), .Y(n2569) );
  OAI2BB1X1 U6312 ( .A0N(n7177), .A1N(N5016), .B0(n2657), .Y(n2652) );
  AND3X2 U6313 ( .A(n2664), .B(n2665), .C(n2662), .Y(n2660) );
  NAND4X1 U6314 ( .A(n2621), .B(n2622), .C(n2623), .D(n2624), .Y(N5146) );
  AOI222XL U6315 ( .A0(N5091), .A1(n2558), .B0(n5572), .B1(n2557), .C0(N5107), 
        .C1(n2555), .Y(n2621) );
  AOI222XL U6316 ( .A0(n5571), .A1(n2556), .B0(N5123), .B1(n2554), .C0(n5572), 
        .C1(n2552), .Y(n2622) );
  AND4X2 U6317 ( .A(n2630), .B(n2631), .C(n2632), .D(n2633), .Y(n2623) );
  AND3X2 U6318 ( .A(n2658), .B(n2659), .C(n2660), .Y(n2657) );
  AND3X2 U6319 ( .A(n2670), .B(n2671), .C(n2672), .Y(n2662) );
  INVX2 U6320 ( .A(n2732), .Y(n7186) );
  OAI2BB1X1 U6321 ( .A0N(N6478), .A1N(n4993), .B0(n6361), .Y(n3210) );
  OR2X1 U6322 ( .A(n6944), .B(n6387), .Y(n6361) );
  OAI2BB1X1 U6323 ( .A0N(N6272), .A1N(n4996), .B0(n6636), .Y(n3486) );
  OR2X1 U6324 ( .A(n4882), .B(n6661), .Y(n6636) );
  NOR3X1 U6325 ( .A(n1313), .B(N5018), .C(n2652), .Y(n2570) );
  NAND4X1 U6326 ( .A(n2639), .B(n2640), .C(n2641), .D(n2642), .Y(N5145) );
  AOI222XL U6327 ( .A0(n5573), .A1(n2555), .B0(N5059), .B1(n2556), .C0(N5059), 
        .C1(n2557), .Y(n2639) );
  AOI222XL U6328 ( .A0(N5059), .A1(n2552), .B0(n5573), .B1(n2553), .C0(n5573), 
        .C1(n2554), .Y(n2640) );
  NOR4BBX1 U6329 ( .AN(n2666), .BN(n2630), .C(n2667), .D(n2668), .Y(n2641) );
  OAI2BB1X1 U6330 ( .A0N(N6190), .A1N(n4994), .B0(n6746), .Y(n3596) );
  OR2X1 U6331 ( .A(n4872), .B(n6771), .Y(n6746) );
  OAI2BB1X1 U6332 ( .A0N(N6353), .A1N(n4999), .B0(n6525), .Y(n3377) );
  OR2X1 U6333 ( .A(n4905), .B(n6549), .Y(n6525) );
  OAI2BB1X1 U6334 ( .A0N(N6435), .A1N(n4992), .B0(n6417), .Y(n3267) );
  OR2X1 U6335 ( .A(n4936), .B(n6441), .Y(n6417) );
  OAI2BB1X1 U6336 ( .A0N(N6313), .A1N(n4997), .B0(n6580), .Y(n3431) );
  OR2X1 U6337 ( .A(n4873), .B(n6605), .Y(n6580) );
  OAI2BB1X1 U6338 ( .A0N(N6395), .A1N(n5000), .B0(n6470), .Y(n3321) );
  OR2X1 U6339 ( .A(n4889), .B(n6495), .Y(n6470) );
  OAI2BB1X1 U6340 ( .A0N(N6189), .A1N(n4994), .B0(n6747), .Y(n3597) );
  OR2X1 U6341 ( .A(n4924), .B(n6771), .Y(n6747) );
  OAI2BB1X1 U6342 ( .A0N(N6271), .A1N(n4996), .B0(n6637), .Y(n3487) );
  OR2X1 U6343 ( .A(n4935), .B(n6661), .Y(n6637) );
  OAI2BB1X1 U6344 ( .A0N(N6312), .A1N(n4997), .B0(n6581), .Y(n3432) );
  OR2X1 U6345 ( .A(n4925), .B(n6605), .Y(n6581) );
  OAI2BB1X1 U6346 ( .A0N(N6477), .A1N(n4993), .B0(n6362), .Y(n3211) );
  OR2X1 U6347 ( .A(n4859), .B(n6387), .Y(n6362) );
  NAND3X1 U6348 ( .A(N5016), .B(n7177), .C(n2657), .Y(n2564) );
  OAI2BB1X1 U6349 ( .A0N(N6394), .A1N(n5000), .B0(n6471), .Y(n3322) );
  OR2X1 U6350 ( .A(n4941), .B(n6495), .Y(n6471) );
  OAI2BB1X1 U6351 ( .A0N(N6476), .A1N(n4993), .B0(n6363), .Y(n3212) );
  OR2X1 U6352 ( .A(n4910), .B(n6387), .Y(n6363) );
  OAI2BB1X1 U6353 ( .A0N(N6186), .A1N(n4994), .B0(n6751), .Y(n3600) );
  OR2X1 U6354 ( .A(n4878), .B(n6771), .Y(n6751) );
  OAI2BB1X1 U6355 ( .A0N(N6185), .A1N(n4994), .B0(n6752), .Y(n3601) );
  OR2X1 U6356 ( .A(n4931), .B(n6771), .Y(n6752) );
  OAI2BB1X1 U6357 ( .A0N(N6432), .A1N(n4992), .B0(n6421), .Y(n3270) );
  OR2X1 U6358 ( .A(n4888), .B(n6441), .Y(n6421) );
  NOR2X1 U6359 ( .A(n2732), .B(n5380), .Y(n2651) );
  NAND2BX1 U6360 ( .AN(n2659), .B(n2660), .Y(n2563) );
  OAI2BB1X1 U6361 ( .A0N(N6391), .A1N(n5000), .B0(n6475), .Y(n3325) );
  OR2X1 U6362 ( .A(n4891), .B(n6495), .Y(n6475) );
  INVX2 U6363 ( .A(n2671), .Y(n7187) );
  OAI2BB1X1 U6364 ( .A0N(N6350), .A1N(n4999), .B0(n6529), .Y(n3380) );
  OR2X1 U6365 ( .A(n4857), .B(n6549), .Y(n6529) );
  NAND3BX1 U6366 ( .AN(n2658), .B(n2660), .C(n2659), .Y(n2565) );
  OAI2BB1X1 U6367 ( .A0N(N6268), .A1N(n4996), .B0(n6641), .Y(n3490) );
  OR2X1 U6368 ( .A(n4885), .B(n6661), .Y(n6641) );
  OAI2BB1X1 U6369 ( .A0N(N6309), .A1N(n4997), .B0(n6585), .Y(n3435) );
  OR2X1 U6370 ( .A(n4879), .B(n6605), .Y(n6585) );
  OAI2BB1X1 U6371 ( .A0N(N6227), .A1N(n4995), .B0(n6696), .Y(n3545) );
  OR2X1 U6372 ( .A(n4866), .B(n6716), .Y(n6696) );
  OAI2BB1X1 U6373 ( .A0N(N6349), .A1N(n4999), .B0(n6530), .Y(n3381) );
  OR2X1 U6374 ( .A(n4909), .B(n6549), .Y(n6530) );
  OAI2BB1X1 U6375 ( .A0N(N6473), .A1N(n4993), .B0(n6367), .Y(n3215) );
  OR2X1 U6376 ( .A(n4861), .B(n6387), .Y(n6367) );
  NOR2X1 U6377 ( .A(n2685), .B(n2671), .Y(n2680) );
  OAI2BB1X1 U6378 ( .A0N(N6226), .A1N(n4995), .B0(n6697), .Y(n3546) );
  OR2X1 U6379 ( .A(n4919), .B(n6716), .Y(n6697) );
  OAI2BB1X1 U6380 ( .A0N(N6308), .A1N(n4997), .B0(n6586), .Y(n3436) );
  OR2X1 U6381 ( .A(n4929), .B(n6605), .Y(n6586) );
  OAI2BB1X1 U6382 ( .A0N(N6390), .A1N(n5000), .B0(n6476), .Y(n3326) );
  OR2X1 U6383 ( .A(n4943), .B(n6495), .Y(n6476) );
  OAI2BB1X1 U6384 ( .A0N(N6431), .A1N(n4992), .B0(n6422), .Y(n3271) );
  OR2X1 U6385 ( .A(n4940), .B(n6441), .Y(n6422) );
  OAI2BB1X1 U6386 ( .A0N(N6472), .A1N(n4993), .B0(n6368), .Y(n3216) );
  OR2X1 U6387 ( .A(n4912), .B(n6387), .Y(n6368) );
  AND3X2 U6388 ( .A(n7187), .B(n2685), .C(n2734), .Y(n2683) );
  AOI2BB2X1 U6389 ( .B0(n5573), .B1(n5572), .A0N(n7311), .A1N(n2733), .Y(n2734) );
  NOR3BX1 U6390 ( .AN(n2662), .B(n7175), .C(n2664), .Y(n2560) );
  OAI2BB1X1 U6391 ( .A0N(N6267), .A1N(n4996), .B0(n6642), .Y(n3491) );
  OR2X1 U6392 ( .A(n4938), .B(n6661), .Y(n6642) );
  NAND2X1 U6393 ( .A(n7187), .B(n2679), .Y(n2676) );
  OAI211X1 U6394 ( .A0(n5380), .A1(n5573), .B0(n5572), .C0(n5379), .Y(n2679)
         );
  NAND2BX1 U6395 ( .AN(n2670), .B(n2672), .Y(n2635) );
  AOI222XL U6396 ( .A0(N5136), .A1(n2552), .B0(N5144), .B1(n2553), .C0(N5128), 
        .C1(n2554), .Y(n2546) );
  OAI222X1 U6397 ( .A0(n7438), .A1(n2635), .B0(n2669), .B1(n7230), .C0(n7445), 
        .C1(n2634), .Y(n2667) );
  NOR2BX1 U6398 ( .AN(n2673), .B(n2674), .Y(n2669) );
  OR2X1 U6399 ( .A(n2814), .B(n5375), .Y(n1585) );
  NAND4X1 U6400 ( .A(n2673), .B(n2638), .C(n2698), .D(n2699), .Y(n2602) );
  AOI211X1 U6401 ( .A0(n2700), .A1(n2701), .B0(n2619), .C0(n7328), .Y(n2699)
         );
  NAND2X1 U6402 ( .A(n2711), .B(n2712), .Y(n2674) );
  AOI222XL U6403 ( .A0(n2710), .A1(n7045), .B0(n7044), .B1(n7013), .C0(n7328), 
        .C1(n7019), .Y(n2711) );
  AOI222XL U6404 ( .A0(n1779), .A1(n7015), .B0(n7014), .B1(n2713), .C0(n2700), 
        .C1(n7325), .Y(n2712) );
  INVX2 U6405 ( .A(n2705), .Y(n7325) );
  NOR3BX1 U6406 ( .AN(n2715), .B(n5373), .C(n7330), .Y(n1827) );
  NAND2X1 U6407 ( .A(n1827), .B(n5375), .Y(n2800) );
  INVX2 U6408 ( .A(n1313), .Y(n7177) );
  OAI2BB1X1 U6409 ( .A0N(N6223), .A1N(n4995), .B0(n6700), .Y(n3549) );
  OR2X1 U6410 ( .A(n4864), .B(n6716), .Y(n6700) );
  NAND2X1 U6411 ( .A(n2715), .B(n7330), .Y(n1743) );
  NOR2X1 U6412 ( .A(n1743), .B(n5375), .Y(n2718) );
  NAND2X1 U6413 ( .A(n5373), .B(n2718), .Y(n2805) );
  OAI211X1 U6414 ( .A0(n2704), .A1(n2705), .B0(n2706), .C0(n2707), .Y(n2637)
         );
  AOI22X1 U6415 ( .A0(n7016), .A1(n7021), .B0(n7046), .B1(n7025), .Y(n2707) );
  AOI33X1 U6416 ( .A0(n7014), .A1(n5376), .A2(n2708), .B0(n7322), .B1(n7035), 
        .B2(n2710), .Y(n2706) );
  INVX2 U6417 ( .A(n2708), .Y(n7322) );
  OR2X1 U6418 ( .A(n7038), .B(n7035), .Y(n2106) );
  INVX2 U6419 ( .A(n5376), .Y(n7035) );
  OAI2BB1X1 U6420 ( .A0N(N6181), .A1N(n4994), .B0(n6756), .Y(n3605) );
  OR2X1 U6421 ( .A(n4926), .B(n6771), .Y(n6756) );
  AOI222XL U6422 ( .A0(N5103), .A1(n2557), .B0(N5135), .B1(n2552), .C0(n5378), 
        .C1(n2556), .Y(n2576) );
  OAI2BB1X1 U6423 ( .A0N(N6428), .A1N(n4992), .B0(n6425), .Y(n3274) );
  OR2X1 U6424 ( .A(n4886), .B(n6441), .Y(n6425) );
  OAI2BB1X1 U6425 ( .A0N(N6387), .A1N(n5000), .B0(n6479), .Y(n3329) );
  OR2X1 U6426 ( .A(n4890), .B(n6495), .Y(n6479) );
  OR2X1 U6427 ( .A(n2814), .B(n7039), .Y(n6552) );
  OAI2BB1X1 U6428 ( .A0N(N6222), .A1N(n4995), .B0(n6701), .Y(n3550) );
  OR2X1 U6429 ( .A(n4915), .B(n6716), .Y(n6701) );
  OAI2BB1X1 U6430 ( .A0N(N6182), .A1N(n4994), .B0(n6755), .Y(n3604) );
  OR2X1 U6431 ( .A(n4875), .B(n6771), .Y(n6755) );
  INVX2 U6432 ( .A(n5374), .Y(n7329) );
  OAI2BB1X1 U6433 ( .A0N(N6264), .A1N(n4996), .B0(n6645), .Y(n3494) );
  OR2X1 U6434 ( .A(n4881), .B(n6661), .Y(n6645) );
  OR2X1 U6435 ( .A(n5376), .B(n7038), .Y(n2788) );
  NAND2X1 U6436 ( .A(n7032), .B(n5374), .Y(n2704) );
  INVX2 U6437 ( .A(n2804), .Y(n7032) );
  AOI222XL U6438 ( .A0(N5112), .A1(n2555), .B0(N5120), .B1(n2556), .C0(N5104), 
        .C1(n2557), .Y(n2545) );
  INVX2 U6439 ( .A(n5377), .Y(N5120) );
  OAI2BB1X1 U6440 ( .A0N(N6386), .A1N(n5000), .B0(n6480), .Y(n3330) );
  OR2X1 U6441 ( .A(n4942), .B(n6495), .Y(n6480) );
  OAI2BB1X1 U6442 ( .A0N(N6427), .A1N(n4992), .B0(n6426), .Y(n3275) );
  OR2X1 U6443 ( .A(n4939), .B(n6441), .Y(n6426) );
  OAI2BB1X1 U6444 ( .A0N(N6305), .A1N(n4997), .B0(n6589), .Y(n3439) );
  OR2X1 U6445 ( .A(n4876), .B(n6605), .Y(n6589) );
  INVX2 U6446 ( .A(n1910), .Y(n7021) );
  OAI2BB1X1 U6447 ( .A0N(N6346), .A1N(n4999), .B0(n6533), .Y(n3384) );
  OR2X1 U6448 ( .A(n4856), .B(n6549), .Y(n6533) );
  XOR2X1 U6449 ( .A(n7038), .B(n5374), .Y(n2708) );
  OR2X1 U6450 ( .A(n5375), .B(n6390), .Y(n1484) );
  OAI2BB1X1 U6451 ( .A0N(N6263), .A1N(n4996), .B0(n6646), .Y(n3495) );
  OR2X1 U6452 ( .A(n4932), .B(n6661), .Y(n6646) );
  OAI2BB1X1 U6453 ( .A0N(N6469), .A1N(n4993), .B0(n6371), .Y(n3219) );
  OR2X1 U6454 ( .A(n4860), .B(n6387), .Y(n6371) );
  OAI2BB1X1 U6455 ( .A0N(N6468), .A1N(n4993), .B0(n6372), .Y(n3220) );
  OR2X1 U6456 ( .A(n4911), .B(n6387), .Y(n6372) );
  OAI2BB1X1 U6457 ( .A0N(N6345), .A1N(n4999), .B0(n6534), .Y(n3385) );
  OR2X1 U6458 ( .A(n4908), .B(n6549), .Y(n6534) );
  OAI2BB1X1 U6459 ( .A0N(N6304), .A1N(n4997), .B0(n6590), .Y(n3440) );
  OR2X1 U6460 ( .A(n4928), .B(n6605), .Y(n6590) );
  NAND2X1 U6461 ( .A(n5375), .B(n2701), .Y(n2696) );
  NOR2X1 U6462 ( .A(n1743), .B(n5373), .Y(n2701) );
  OR2X1 U6463 ( .A(n5374), .B(n2696), .Y(n6777) );
  AOI221XL U6464 ( .A0(n2701), .A1(n7320), .B0(n7045), .B1(n7044), .C0(n2722), 
        .Y(n2673) );
  OAI32X1 U6465 ( .A0(n7039), .A1(n1743), .A2(n2723), .B0(n7038), .B1(n2698), 
        .Y(n2722) );
  INVX2 U6466 ( .A(n2814), .Y(n7046) );
  INVX2 U6467 ( .A(n5375), .Y(n7039) );
  INVX2 U6468 ( .A(n2665), .Y(n7175) );
  NOR2X1 U6469 ( .A(n2804), .B(n5374), .Y(n1779) );
  AOI22X1 U6470 ( .A0(N5111), .A1(n2555), .B0(N5095), .B1(n2558), .Y(n2575) );
  INVX2 U6471 ( .A(n5373), .Y(n7040) );
  NAND2X1 U6472 ( .A(n7327), .B(n5374), .Y(n2689) );
  NAND2X1 U6473 ( .A(n7034), .B(n2692), .Y(n2630) );
  OAI31X1 U6474 ( .A0(n1863), .A1(n5374), .A2(n7025), .B0(n2108), .Y(n2692) );
  AOI22X1 U6475 ( .A0(N5096), .A1(n2558), .B0(N5072), .B1(n2559), .Y(n2544) );
  OAI2BB1X1 U6476 ( .A0N(N6260), .A1N(n4996), .B0(n6649), .Y(n3498) );
  OR2X1 U6477 ( .A(n4871), .B(n6661), .Y(n6649) );
  AND2X1 U6478 ( .A(n2785), .B(n2786), .Y(n2784) );
  NOR4BBX1 U6479 ( .AN(n2757), .BN(n2756), .C(n2787), .D(n7205), .Y(n2786) );
  NOR4X1 U6480 ( .A(n2795), .B(n2748), .C(n2539), .D(n2754), .Y(n2785) );
  NAND4X1 U6481 ( .A(n2686), .B(n2765), .C(n2601), .D(n2777), .Y(n2787) );
  NAND2BX1 U6482 ( .AN(n5373), .B(n2718), .Y(n6775) );
  OR2X1 U6483 ( .A(n96), .B(n5442), .Y(n7230) );
  INVX2 U6484 ( .A(n7232), .Y(n5434) );
  NAND2X1 U6485 ( .A(n2784), .B(n117), .Y(n2735) );
  OAI2BB1X1 U6486 ( .A0N(N6424), .A1N(n4992), .B0(n6429), .Y(n3278) );
  OR2X1 U6487 ( .A(n4874), .B(n6441), .Y(n6429) );
  NOR3BX1 U6488 ( .AN(n1312), .B(n1313), .C(n1314), .Y(n1269) );
  AND2X1 U6489 ( .A(n1269), .B(n5570), .Y(n1237) );
  NAND3X1 U6490 ( .A(n5572), .B(n5569), .C(n1237), .Y(n1233) );
  OAI2BB2X1 U6491 ( .B0(n1281), .B1(n7478), .A0N(N4934), .A1N(n7181), .Y(n3151) );
  OAI2BB2X1 U6492 ( .B0(n1281), .B1(n7477), .A0N(N4933), .A1N(n7181), .Y(n3152) );
  OAI2BB2X1 U6493 ( .B0(n1281), .B1(n7476), .A0N(N4932), .A1N(n7181), .Y(n3153) );
  NAND3X1 U6494 ( .A(n1237), .B(n5572), .C(n5568), .Y(n1280) );
  NAND3X1 U6495 ( .A(n1237), .B(n5569), .C(n5571), .Y(n1247) );
  OAI2BB2X1 U6496 ( .B0(n1271), .B1(n7471), .A0N(N4917), .A1N(n7182), .Y(n3144) );
  OAI2BB2X1 U6497 ( .B0(n1271), .B1(n7470), .A0N(N4916), .A1N(n7182), .Y(n3145) );
  OAI2BB2X1 U6498 ( .B0(n1271), .B1(n7469), .A0N(N4915), .A1N(n7182), .Y(n3146) );
  NOR3BX1 U6499 ( .AN(n1269), .B(n5571), .C(n5570), .Y(n1258) );
  NAND2X1 U6500 ( .A(n1258), .B(n5569), .Y(n1257) );
  OAI2BB1X1 U6501 ( .A0N(N6219), .A1N(n4995), .B0(n6704), .Y(n3553) );
  OR2X1 U6502 ( .A(n4862), .B(n6716), .Y(n6704) );
  OR2X1 U6503 ( .A(n96), .B(n5464), .Y(n7206) );
  INVX2 U6504 ( .A(n111), .Y(n5467) );
  OAI2BB1X1 U6505 ( .A0N(N6178), .A1N(n4994), .B0(n6759), .Y(n3608) );
  OR2X1 U6506 ( .A(n4867), .B(n6771), .Y(n6759) );
  OAI2BB1X1 U6507 ( .A0N(N6342), .A1N(n4999), .B0(n6537), .Y(n3388) );
  OR2X1 U6508 ( .A(n4852), .B(n6549), .Y(n6537) );
  OAI2BB1X1 U6509 ( .A0N(N6465), .A1N(n4993), .B0(n6375), .Y(n3223) );
  OR2X1 U6510 ( .A(n4855), .B(n6387), .Y(n6375) );
  INVX2 U6511 ( .A(n2783), .Y(n7028) );
  OAI2BB1X1 U6512 ( .A0N(N6259), .A1N(n4996), .B0(n6650), .Y(n3499) );
  OR2X1 U6513 ( .A(n4923), .B(n6661), .Y(n6650) );
  OAI2BB1X1 U6514 ( .A0N(N6218), .A1N(n4995), .B0(n6705), .Y(n3554) );
  OR2X1 U6515 ( .A(n4914), .B(n6716), .Y(n6705) );
  OAI2BB1X1 U6516 ( .A0N(N6383), .A1N(n5000), .B0(n6483), .Y(n3333) );
  OR2X1 U6517 ( .A(n4883), .B(n6495), .Y(n6483) );
  OAI2BB1X1 U6518 ( .A0N(N6301), .A1N(n4997), .B0(n6593), .Y(n3443) );
  OR2X1 U6519 ( .A(n4868), .B(n6605), .Y(n6593) );
  XOR2X1 U6520 ( .A(n5376), .B(n5374), .Y(n2717) );
  OAI2BB1X1 U6521 ( .A0N(N6177), .A1N(n4994), .B0(n6760), .Y(n3609) );
  OR2X1 U6522 ( .A(n4917), .B(n6771), .Y(n6760) );
  OAI2BB1X1 U6523 ( .A0N(N6341), .A1N(n4999), .B0(n6538), .Y(n3389) );
  OR2X1 U6524 ( .A(n4904), .B(n6549), .Y(n6538) );
  OAI2BB1X1 U6525 ( .A0N(N6382), .A1N(n5000), .B0(n6484), .Y(n3334) );
  OR2X1 U6526 ( .A(n4937), .B(n6495), .Y(n6484) );
  OAI2BB1X1 U6527 ( .A0N(N6300), .A1N(n4997), .B0(n6594), .Y(n3444) );
  OR2X1 U6528 ( .A(n4921), .B(n6605), .Y(n6594) );
  OAI2BB1X1 U6529 ( .A0N(N6464), .A1N(n4993), .B0(n6376), .Y(n3224) );
  OR2X1 U6530 ( .A(n4907), .B(n6387), .Y(n6376) );
  OAI2BB1X1 U6531 ( .A0N(N6423), .A1N(n4992), .B0(n6430), .Y(n3279) );
  OR2X1 U6532 ( .A(n4930), .B(n6441), .Y(n6430) );
  NAND3X1 U6533 ( .A(n1269), .B(n5569), .C(n1270), .Y(n1268) );
  OAI2BB2X1 U6534 ( .B0(n1259), .B1(n7464), .A0N(N4900), .A1N(n7185), .Y(n3137) );
  OAI2BB2X1 U6535 ( .B0(n1259), .B1(n7463), .A0N(N4899), .A1N(n7185), .Y(n3138) );
  OAI2BB2X1 U6536 ( .B0(n1259), .B1(n7462), .A0N(N4898), .A1N(n7185), .Y(n3139) );
  NAND4X1 U6537 ( .A(n2768), .B(n2778), .C(n2779), .D(n2780), .Y(N4778) );
  NOR4BX1 U6538 ( .AN(n2774), .B(n2781), .C(n7205), .D(n7028), .Y(n2780) );
  NAND2X1 U6539 ( .A(n7190), .B(n5379), .Y(n2778) );
  AOI22X1 U6540 ( .A0(n2739), .A1(n5571), .B0(n2737), .B1(N5059), .Y(n2779) );
  NOR2X1 U6541 ( .A(n7168), .B(n102), .Y(n2376) );
  OAI2BB2X1 U6542 ( .B0(n7304), .B1(n4848), .A0N(N4586), .A1N(n2376), .Y(n4024) );
  OAI2BB2X1 U6543 ( .B0(n7302), .B1(n4848), .A0N(N4585), .A1N(n2376), .Y(n4026) );
  OAI2BB2X1 U6544 ( .B0(n7305), .B1(n4848), .A0N(N4587), .A1N(n2376), .Y(n4023) );
  OAI2BB2X1 U6545 ( .B0(n7313), .B1(n4848), .A0N(N4597), .A1N(n2376), .Y(n4013) );
  OAI2BB2X1 U6546 ( .B0(N5120), .B1(n4848), .A0N(N4596), .A1N(n2376), .Y(n4014) );
  OAI2BB2X1 U6547 ( .B0(n5567), .B1(n4848), .A0N(N4594), .A1N(n2376), .Y(n4016) );
  OAI2BB2X1 U6548 ( .B0(n5569), .B1(n4848), .A0N(N4593), .A1N(n2376), .Y(n4017) );
  OAI2BB2X1 U6549 ( .B0(n5570), .B1(n4848), .A0N(N4592), .A1N(n2376), .Y(n4018) );
  OAI2BB2X1 U6550 ( .B0(n5572), .B1(n4848), .A0N(N4591), .A1N(n2376), .Y(n4019) );
  OR2X1 U6551 ( .A(n5415), .B(n96), .Y(n6776) );
  OAI2BB2X1 U6552 ( .B0(n4848), .B1(n5573), .A0N(N4590), .A1N(n2376), .Y(n4020) );
  INVX2 U6553 ( .A(n2539), .Y(n7189) );
  NAND2X1 U6554 ( .A(n7203), .B(n2362), .Y(n2354) );
  OAI2BB1X1 U6555 ( .A0N(N4695), .A1N(n7042), .B0(n5896), .Y(n4000) );
  OR2X1 U6556 ( .A(n2354), .B(n7035), .Y(n5896) );
  OAI2BB2X1 U6557 ( .B0(n7331), .B1(n2354), .A0N(N4700), .A1N(n7042), .Y(n3994) );
  OAI2BB2X1 U6558 ( .B0(n7330), .B1(n2354), .A0N(N4698), .A1N(n7042), .Y(n3996) );
  NOR2X1 U6559 ( .A(n1910), .B(n7329), .Y(n1561) );
  INVX2 U6560 ( .A(n132), .Y(n7170) );
  INVX2 U6561 ( .A(N7651), .Y(n5253) );
  OAI2BB2X1 U6562 ( .B0(N7652), .B1(n5252), .A0N(n5007), .A1N(N7652), .Y(N9857) );
  OR2X1 U6563 ( .A(n5217), .B(n5216), .Y(n5007) );
  NAND3X1 U6564 ( .A(n7004), .B(n6998), .C(n6997), .Y(n6999) );
  INVX2 U6565 ( .A(n6993), .Y(n6998) );
  NOR2BX1 U6566 ( .AN(n7290), .B(n168), .Y(n6996) );
  INVX2 U6567 ( .A(n7070), .Y(n7072) );
  OAI221X1 U6568 ( .A0(n584), .A1(n7576), .B0(n586), .B1(N7799), .C0(n588), 
        .Y(n583) );
  OAI221X1 U6569 ( .A0(n192), .A1(n193), .B0(n194), .B1(n7243), .C0(n196), .Y(
        n165) );
  NAND4X1 U6570 ( .A(n274), .B(n275), .C(n276), .D(n277), .Y(n164) );
  INVX2 U6571 ( .A(N7610), .Y(n5208) );
  OAI2BB2X1 U6572 ( .B0(N7611), .B1(n5207), .A0N(n5008), .A1N(N7611), .Y(N9808) );
  OR2X1 U6573 ( .A(n5172), .B(n5171), .Y(n5008) );
  INVX2 U6574 ( .A(n7065), .Y(n7067) );
  INVX2 U6575 ( .A(n2362), .Y(n7042) );
  INVX2 U6576 ( .A(N7692), .Y(n5298) );
  OAI2BB2X1 U6577 ( .B0(N7693), .B1(n5297), .A0N(n5009), .A1N(N7693), .Y(N9906) );
  OR2X1 U6578 ( .A(n5262), .B(n5261), .Y(n5009) );
  INVX2 U6579 ( .A(n7075), .Y(n7077) );
  OAI2BB1X1 U6580 ( .A0N(N6174), .A1N(n4994), .B0(n6765), .Y(n3612) );
  OR2X1 U6581 ( .A(n4869), .B(n6771), .Y(n6765) );
  OAI2BB1X1 U6582 ( .A0N(N6215), .A1N(n4995), .B0(n6710), .Y(n3557) );
  OR2X1 U6583 ( .A(n4863), .B(n6716), .Y(n6710) );
  NOR2X1 U6584 ( .A(n2689), .B(n1910), .Y(n2072) );
  OAI2BB1X1 U6585 ( .A0N(N6379), .A1N(n5000), .B0(n6489), .Y(n3337) );
  OR2X1 U6586 ( .A(n4887), .B(n6495), .Y(n6489) );
  OAI2BB1X1 U6587 ( .A0N(N6256), .A1N(n4996), .B0(n6655), .Y(n3502) );
  OR2X1 U6588 ( .A(n4877), .B(n6661), .Y(n6655) );
  INVX2 U6589 ( .A(N7650), .Y(n5254) );
  NAND2X1 U6590 ( .A(N7980), .B(n4952), .Y(n295) );
  OAI2BB1X1 U6591 ( .A0N(N6420), .A1N(n4992), .B0(n6435), .Y(n3282) );
  OR2X1 U6592 ( .A(n4880), .B(n6441), .Y(n6435) );
  INVX2 U6593 ( .A(n2531), .Y(n5897) );
  AOI222XL U6594 ( .A0(n464), .A1(n792), .B0(n349), .B1(n793), .C0(n346), .C1(
        n794), .Y(n791) );
  NAND4X1 U6595 ( .A(n7582), .B(n7583), .C(N7799), .D(n801), .Y(n792) );
  NAND4X1 U6596 ( .A(n7563), .B(n7564), .C(N7871), .D(n799), .Y(n793) );
  NAND4X1 U6597 ( .A(n7591), .B(n7592), .C(n4902), .D(n797), .Y(n794) );
  AOI222XL U6598 ( .A0(n780), .A1(n117), .B0(n7005), .B1(n5466), .C0(n782), 
        .C1(n7004), .Y(n7006) );
  NAND4X1 U6599 ( .A(n739), .B(n873), .C(n874), .D(n875), .Y(n780) );
  OR4X2 U6600 ( .A(n784), .B(n785), .C(n786), .D(n787), .Y(n782) );
  NAND4X1 U6601 ( .A(n823), .B(n862), .C(n739), .D(n863), .Y(n777) );
  AOI211X1 U6602 ( .A0(n7264), .A1(n7250), .B0(n865), .C0(n812), .Y(n863) );
  OAI22X1 U6603 ( .A0(n861), .A1(n745), .B0(n7251), .B1(n867), .Y(n865) );
  AND2X1 U6604 ( .A(n925), .B(n923), .Y(n929) );
  NAND2X1 U6605 ( .A(n283), .B(n190), .Y(n918) );
  INVX2 U6606 ( .A(N7609), .Y(n5209) );
  NAND2X1 U6607 ( .A(n7259), .B(n7529), .Y(n928) );
  INVX2 U6608 ( .A(n188), .Y(n7257) );
  NAND4BX1 U6609 ( .AN(n821), .B(n822), .C(n823), .D(n824), .Y(n784) );
  AOI221XL U6610 ( .A0(n466), .A1(n825), .B0(n600), .B1(n826), .C0(n827), .Y(
        n824) );
  NAND4X1 U6611 ( .A(n4901), .B(n7546), .C(N7943), .D(n846), .Y(n826) );
  NAND4X1 U6612 ( .A(n7600), .B(n7601), .C(N7727), .D(n849), .Y(n825) );
  NOR2X1 U6613 ( .A(n190), .B(n171), .Y(n715) );
  NOR2X1 U6614 ( .A(n188), .B(n171), .Y(n590) );
  NOR2X1 U6615 ( .A(n5363), .B(n800), .Y(n349) );
  OAI2BB1X1 U6616 ( .A0N(N6338), .A1N(n4999), .B0(n6543), .Y(n3392) );
  OR2X1 U6617 ( .A(n4853), .B(n6549), .Y(n6543) );
  OAI2BB1X1 U6618 ( .A0N(N6297), .A1N(n4997), .B0(n6599), .Y(n3447) );
  OR2X1 U6619 ( .A(n4870), .B(n6605), .Y(n6599) );
  OAI2BB1X1 U6620 ( .A0N(N6461), .A1N(n4993), .B0(n6381), .Y(n3227) );
  OR2X1 U6621 ( .A(n4858), .B(n6387), .Y(n6381) );
  OAI22X1 U6622 ( .A0(n297), .A1(n4912), .B0(n295), .B1(n4861), .Y(n313) );
  INVX2 U6623 ( .A(N7691), .Y(n5299) );
  OAI2BB2X1 U6624 ( .B0(N7526), .B1(n5117), .A0N(n5010), .A1N(N7526), .Y(N9710) );
  OR2X1 U6625 ( .A(n5082), .B(n5081), .Y(n5010) );
  INVX2 U6626 ( .A(N7525), .Y(n5118) );
  INVX2 U6627 ( .A(n7055), .Y(n7057) );
  INVX2 U6628 ( .A(N7524), .Y(n5119) );
  OAI22X1 U6629 ( .A0(n7170), .A1(n7036), .B0(n132), .B1(n7193), .Y(n2852) );
  AOI2BB2X1 U6630 ( .B0(n6986), .B1(n117), .A0N(n5464), .A1N(n6985), .Y(n7001)
         );
  OR2X1 U6631 ( .A(n732), .B(n733), .Y(n6986) );
  AOI221XL U6632 ( .A0(n743), .A1(n7041), .B0(n742), .B1(n6984), .C0(n722), 
        .Y(n6985) );
  OAI32X1 U6633 ( .A0(n734), .A1(n7285), .A2(n7261), .B0(n737), .B1(n7245), 
        .Y(n733) );
  INVX2 U6634 ( .A(n7050), .Y(n7052) );
  AND2X1 U6635 ( .A(N9661), .B(n7285), .Y(n197) );
  INVX2 U6636 ( .A(N7480), .Y(n5073) );
  NOR2X1 U6637 ( .A(n4952), .B(N7980), .Y(n301) );
  NAND2X1 U6638 ( .A(n858), .B(n859), .Y(n815) );
  NOR4BBX1 U6639 ( .AN(n586), .BN(n584), .C(n726), .D(n725), .Y(n859) );
  AOI221XL U6640 ( .A0(n199), .A1(n860), .B0(n7279), .B1(n7249), .C0(n345), 
        .Y(n858) );
  NAND2X1 U6641 ( .A(n861), .B(n5362), .Y(n860) );
  NOR2X1 U6642 ( .A(n7192), .B(n2539), .Y(N5258) );
  NAND2X1 U6643 ( .A(N7872), .B(N7871), .Y(n359) );
  NAND2X1 U6644 ( .A(N7764), .B(n4902), .Y(n416) );
  NOR2X1 U6645 ( .A(n283), .B(n171), .Y(n714) );
  NOR2X1 U6646 ( .A(n5363), .B(n171), .Y(n466) );
  NAND2X1 U6647 ( .A(n2524), .B(n2531), .Y(n884) );
  NOR3BX1 U6648 ( .AN(n2525), .B(n7292), .C(n4849), .Y(n2422) );
  NAND2X1 U6649 ( .A(n2493), .B(n2422), .Y(n178) );
  OAI22X1 U6650 ( .A0(n297), .A1(n4910), .B0(n295), .B1(n4859), .Y(n328) );
  INVX2 U6651 ( .A(n297), .Y(n6947) );
  OAI2BB2X1 U6652 ( .B0(N7570), .B1(n5162), .A0N(n5011), .A1N(N7570), .Y(N9759) );
  OR2X1 U6653 ( .A(n5127), .B(n5126), .Y(n5011) );
  INVX2 U6654 ( .A(N7569), .Y(n5163) );
  INVX2 U6655 ( .A(n7060), .Y(n7062) );
  OAI2BB1X1 U6656 ( .A0N(N6214), .A1N(n4995), .B0(n6711), .Y(n3558) );
  OR2X1 U6657 ( .A(n4913), .B(n6716), .Y(n6711) );
  NAND2X1 U6658 ( .A(n2526), .B(n2524), .Y(n182) );
  OAI2BB1X1 U6659 ( .A0N(N6173), .A1N(n4994), .B0(n6766), .Y(n3613) );
  OR2X1 U6660 ( .A(n4918), .B(n6771), .Y(n6766) );
  NAND2X1 U6661 ( .A(n2526), .B(n2493), .Y(n272) );
  OAI22X1 U6662 ( .A0(n361), .A1(n4909), .B0(n359), .B1(n4857), .Y(n377) );
  OAI2BB1X1 U6663 ( .A0N(N6419), .A1N(n4992), .B0(n6436), .Y(n3283) );
  OR2X1 U6664 ( .A(n4927), .B(n6441), .Y(n6436) );
  OAI22X1 U6665 ( .A0(n418), .A1(n4919), .B0(n416), .B1(n4866), .Y(n434) );
  NOR2X1 U6666 ( .A(n7168), .B(n7192), .Y(N5387) );
  NAND2X1 U6667 ( .A(n2520), .B(n2531), .Y(n882) );
  INVX2 U6668 ( .A(N7648), .Y(n5256) );
  INVX2 U6669 ( .A(n800), .Y(n7272) );
  NOR2X1 U6670 ( .A(n190), .B(n182), .Y(n345) );
  AND2X1 U6671 ( .A(n2520), .B(n2526), .Y(n199) );
  NAND2X1 U6672 ( .A(n2493), .B(n2531), .Y(n867) );
  INVX2 U6673 ( .A(n300), .Y(n6960) );
  NAND2X1 U6674 ( .A(n2524), .B(n7291), .Y(n761) );
  INVX2 U6675 ( .A(N7981), .Y(n7534) );
  INVX2 U6676 ( .A(N7607), .Y(n5211) );
  INVX2 U6677 ( .A(n5361), .Y(n7255) );
  NAND2X1 U6678 ( .A(n5362), .B(n193), .Y(n857) );
  NAND2X1 U6679 ( .A(n7251), .B(n5361), .Y(n870) );
  OAI2BB1X1 U6680 ( .A0N(N6296), .A1N(n4997), .B0(n6600), .Y(n3448) );
  OR2X1 U6681 ( .A(n4920), .B(n6605), .Y(n6600) );
  NOR2X1 U6682 ( .A(n4902), .B(N7764), .Y(n422) );
  INVX2 U6683 ( .A(n7110), .Y(n7111) );
  INVX2 U6684 ( .A(N7478), .Y(n5074) );
  NOR2X1 U6685 ( .A(N7871), .B(N7872), .Y(n365) );
  NOR2X1 U6686 ( .A(n188), .B(n182), .Y(n725) );
  NOR2X1 U6687 ( .A(n5361), .B(n182), .Y(n726) );
  NOR2X1 U6688 ( .A(n283), .B(n178), .Y(n721) );
  OAI2BB1X1 U6689 ( .A0N(N6337), .A1N(n4999), .B0(n6544), .Y(n3393) );
  OR2X1 U6690 ( .A(n4903), .B(n6549), .Y(n6544) );
  INVX2 U6691 ( .A(N7689), .Y(n5301) );
  NAND3X1 U6692 ( .A(n7292), .B(n4849), .C(n2525), .Y(n2494) );
  INVX2 U6693 ( .A(n745), .Y(n7275) );
  OAI2BB1X1 U6694 ( .A0N(N6378), .A1N(n5000), .B0(n6490), .Y(n3338) );
  OR2X1 U6695 ( .A(n4933), .B(n6495), .Y(n6490) );
  OAI2BB1X1 U6696 ( .A0N(N6460), .A1N(n4993), .B0(n6382), .Y(n3228) );
  OR2X1 U6697 ( .A(n4906), .B(n6387), .Y(n6382) );
  OAI2BB1X1 U6698 ( .A0N(N6255), .A1N(n4996), .B0(n6656), .Y(n3503) );
  OR2X1 U6699 ( .A(n4922), .B(n6661), .Y(n6656) );
  NAND2X1 U6700 ( .A(n2520), .B(n7291), .Y(n802) );
  OAI22X1 U6701 ( .A0(n361), .A1(n4905), .B0(n359), .B1(n4854), .Y(n392) );
  INVX2 U6702 ( .A(n361), .Y(n6923) );
  OAI22X1 U6703 ( .A0(n418), .A1(n4916), .B0(n416), .B1(n4865), .Y(n449) );
  INVX2 U6704 ( .A(n418), .Y(n6899) );
  INVX2 U6705 ( .A(N7568), .Y(n5164) );
  NAND2X1 U6706 ( .A(N7944), .B(N7943), .Y(n610) );
  NOR2X1 U6707 ( .A(n761), .B(n5362), .Y(n764) );
  NOR2X1 U6708 ( .A(n272), .B(n5361), .Y(n589) );
  NOR2X1 U6709 ( .A(n761), .B(n193), .Y(n765) );
  NOR2X1 U6710 ( .A(n5362), .B(n272), .Y(n591) );
  INVX2 U6711 ( .A(n421), .Y(n6912) );
  INVX2 U6712 ( .A(n364), .Y(n6936) );
  INVX2 U6713 ( .A(N7873), .Y(n7560) );
  INVX2 U6714 ( .A(N7765), .Y(n7588) );
  OAI22X1 U6715 ( .A0(n612), .A1(n4940), .B0(n610), .B1(n4888), .Y(n628) );
  INVX2 U6716 ( .A(N7982), .Y(n7535) );
  AOI22X1 U6717 ( .A0(n464), .A1(n465), .B0(n466), .B1(n467), .Y(n274) );
  OAI222X1 U6718 ( .A0(n468), .A1(n7599), .B0(N7731), .B1(n470), .C0(n471), 
        .C1(n5026), .Y(n467) );
  OAI222X1 U6719 ( .A0(n524), .A1(n7581), .B0(N7803), .B1(n526), .C0(n527), 
        .C1(n5028), .Y(n465) );
  AOI22X1 U6720 ( .A0(n473), .A1(n7597), .B0(N7729), .B1(n475), .Y(n471) );
  INVX2 U6721 ( .A(n7085), .Y(n7086) );
  INVX2 U6722 ( .A(n7098), .Y(n7099) );
  NAND2X1 U6723 ( .A(N7800), .B(N7799), .Y(n532) );
  NAND2X1 U6724 ( .A(N7728), .B(N7727), .Y(n476) );
  INVX2 U6725 ( .A(n283), .Y(n7244) );
  INVX2 U6726 ( .A(n190), .Y(n7260) );
  NAND4X1 U6727 ( .A(n882), .B(n745), .C(n884), .D(n896), .Y(n840) );
  NOR2X1 U6728 ( .A(n7277), .B(n7261), .Y(n896) );
  NAND2X1 U6729 ( .A(N7836), .B(N7835), .Y(n229) );
  NAND2X1 U6730 ( .A(N7836), .B(n5364), .Y(n227) );
  INVX2 U6731 ( .A(N7522), .Y(n5121) );
  NAND2X1 U6732 ( .A(N7908), .B(n5365), .Y(n668) );
  NOR2X1 U6733 ( .A(N7943), .B(N7944), .Y(n616) );
  NAND2X1 U6734 ( .A(n2520), .B(n2422), .Y(n169) );
  NOR2X1 U6735 ( .A(n169), .B(n193), .Y(n720) );
  NAND2X1 U6736 ( .A(n2524), .B(n2422), .Y(n831) );
  NOR2X1 U6737 ( .A(n169), .B(n5361), .Y(n718) );
  NAND2X1 U6738 ( .A(N7908), .B(N7907), .Y(n666) );
  OAI22X1 U6739 ( .A0(n534), .A1(n4938), .B0(n532), .B1(n4885), .Y(n550) );
  OAI22X1 U6740 ( .A0(n478), .A1(n4931), .B0(n476), .B1(n4878), .Y(n494) );
  NOR2X1 U6741 ( .A(n831), .B(n190), .Y(n719) );
  INVX2 U6742 ( .A(N7476), .Y(n5076) );
  OAI22X1 U6743 ( .A0(n227), .A1(n4929), .B0(n229), .B1(n4879), .Y(n231) );
  NOR2X1 U6744 ( .A(N7835), .B(N7836), .Y(n225) );
  OAI22X1 U6745 ( .A0(n668), .A1(n4943), .B0(n666), .B1(n4891), .Y(n684) );
  OAI22X1 U6746 ( .A0(n612), .A1(n4936), .B0(n610), .B1(n4884), .Y(n643) );
  NOR2X1 U6747 ( .A(n831), .B(n283), .Y(n344) );
  INVX2 U6748 ( .A(n612), .Y(n6827) );
  NOR2X1 U6749 ( .A(N7907), .B(N7908), .Y(n672) );
  NOR2X1 U6750 ( .A(n5364), .B(N7836), .Y(n224) );
  NOR2X1 U6751 ( .A(N7799), .B(N7800), .Y(n538) );
  NOR2X1 U6752 ( .A(N7727), .B(N7728), .Y(n482) );
  INVX2 U6753 ( .A(N7766), .Y(n7589) );
  INVX2 U6754 ( .A(N7874), .Y(n7561) );
  INVX2 U6755 ( .A(N7566), .Y(n5166) );
  NOR2X1 U6756 ( .A(n831), .B(n5362), .Y(n597) );
  INVX2 U6757 ( .A(n193), .Y(n7249) );
  INVX2 U6758 ( .A(n7093), .Y(n7095) );
  INVX2 U6759 ( .A(N7840), .Y(n7571) );
  NOR2X1 U6760 ( .A(n5365), .B(N7908), .Y(n671) );
  INVX2 U6761 ( .A(n615), .Y(n6840) );
  NOR4X1 U6762 ( .A(n7305), .B(n7304), .C(n7302), .D(n7303), .Y(n1312) );
  INVX2 U6763 ( .A(N7945), .Y(n7543) );
  INVX2 U6764 ( .A(n7106), .Y(n7107) );
  OAI22X1 U6765 ( .A0(n534), .A1(n4935), .B0(n532), .B1(n4882), .Y(n565) );
  OAI22X1 U6766 ( .A0(n478), .A1(n4924), .B0(n476), .B1(n4872), .Y(n509) );
  INVX2 U6767 ( .A(n534), .Y(n6851) );
  INVX2 U6768 ( .A(n478), .Y(n6875) );
  OAI22X1 U6769 ( .A0(n227), .A1(n4925), .B0(n229), .B1(n4873), .Y(n246) );
  NAND2X1 U6770 ( .A(N9425), .B(N7419), .Y(n734) );
  INVX2 U6771 ( .A(N7432), .Y(n5346) );
  OAI22X1 U6772 ( .A0(n668), .A1(n4941), .B0(n666), .B1(n4889), .Y(n699) );
  INVX2 U6773 ( .A(n537), .Y(n6864) );
  INVX2 U6774 ( .A(n481), .Y(n6888) );
  INVX2 U6775 ( .A(N7801), .Y(n7579) );
  INVX2 U6776 ( .A(N7729), .Y(n7597) );
  INVX2 U6777 ( .A(n7102), .Y(n7103) );
  INVX2 U6778 ( .A(N7837), .Y(n7569) );
  INVX2 U6779 ( .A(n7080), .Y(n7082) );
  INVX2 U6780 ( .A(N7479), .Y(n5072) );
  INVX2 U6781 ( .A(n5379), .Y(n7311) );
  INVX2 U6782 ( .A(n7089), .Y(n7090) );
  INVX2 U6783 ( .A(N7909), .Y(n7551) );
  OAI211X1 U6784 ( .A0(n744), .A1(n745), .B0(n7240), .C0(n747), .Y(n722) );
  AND2X1 U6785 ( .A(n771), .B(n772), .Y(n744) );
  INVX2 U6786 ( .A(n732), .Y(n7240) );
  AOI222XL U6787 ( .A0(n7286), .A1(n749), .B0(n7264), .B1(n751), .C0(n7277), 
        .C1(n753), .Y(n747) );
  INVX2 U6788 ( .A(N7649), .Y(n5255) );
  INVX2 U6789 ( .A(N7983), .Y(n7536) );
  INVX2 U6790 ( .A(n111), .Y(n5465) );
  INVX2 U6791 ( .A(N7946), .Y(n7544) );
  INVX2 U6792 ( .A(n5380), .Y(n7310) );
  INVX2 U6793 ( .A(N7608), .Y(n5210) );
  INVX2 U6794 ( .A(N7838), .Y(n7570) );
  OAI22X1 U6795 ( .A0(n6977), .A1(n6966), .B0(n6975), .B1(n6965), .Y(n6967) );
  NOR2X1 U6796 ( .A(n117), .B(n5895), .Y(n5012) );
  INVX2 U6797 ( .A(n5012), .Y(n7007) );
  INVX2 U6798 ( .A(n7232), .Y(n5435) );
  INVX2 U6799 ( .A(N7690), .Y(n5300) );
  INVX2 U6800 ( .A(N7910), .Y(n7552) );
  INVX2 U6801 ( .A(N7730), .Y(n7598) );
  INVX2 U6802 ( .A(N7802), .Y(n7580) );
  INVX2 U6803 ( .A(n2422), .Y(n5899) );
  BUFX2 U6804 ( .A(n140), .Y(n5350) );
  OAI2BB1X1 U6805 ( .A0N(n7034), .A1N(n5015), .B0(n5902), .Y(n140) );
  OAI2BB1X1 U6806 ( .A0N(n6791), .A1N(n5901), .B0(n5900), .Y(n5902) );
  INVX2 U6807 ( .A(n5362), .Y(n7254) );
  INVX2 U6808 ( .A(N7430), .Y(n5345) );
  NAND2X1 U6809 ( .A(n7030), .B(n2797), .Y(n2774) );
  NAND4BBX1 U6810 ( .AN(n1944), .BN(n7022), .C(n2798), .D(n2799), .Y(n2797) );
  NAND3X1 U6811 ( .A(n2717), .B(n7038), .C(n7014), .Y(n2798) );
  AOI222XL U6812 ( .A0(n7326), .A1(n7032), .B0(n7044), .B1(n7025), .C0(n7324), 
        .C1(n7013), .Y(n2799) );
  INVX2 U6813 ( .A(N7523), .Y(n5120) );
  NAND3X1 U6814 ( .A(n877), .B(n862), .C(n919), .Y(n818) );
  AOI222XL U6815 ( .A0(n7255), .A1(n7275), .B0(n7264), .B1(n920), .C0(n7277), 
        .C1(n7249), .Y(n919) );
  NAND3X1 U6816 ( .A(n5361), .B(n5362), .C(n188), .Y(n920) );
  INVX2 U6817 ( .A(N7767), .Y(n7590) );
  INVX2 U6818 ( .A(N7875), .Y(n7562) );
  NAND2X1 U6819 ( .A(n7030), .B(n2813), .Y(n2796) );
  OAI221X1 U6820 ( .A0(n1864), .A1(n2814), .B0(n2793), .B1(n1863), .C0(n2815), 
        .Y(n2813) );
  AOI222XL U6821 ( .A0(n7014), .A1(n7045), .B0(n1779), .B1(n7015), .C0(n7044), 
        .C1(n7023), .Y(n2815) );
  NAND2X1 U6822 ( .A(n7030), .B(n2803), .Y(n2762) );
  OAI221X1 U6823 ( .A0(n2804), .A1(n2805), .B0(n2788), .B1(n2689), .C0(n2806), 
        .Y(n2803) );
  AOI221XL U6824 ( .A0(n7043), .A1(n7014), .B0(n2716), .B1(n7324), .C0(n7015), 
        .Y(n2806) );
  NAND2X1 U6825 ( .A(n7030), .B(n2775), .Y(n2807) );
  XOR2X1 U6826 ( .A(n5380), .B(N5059), .Y(n2685) );
  OAI221X1 U6827 ( .A0(N7688), .A1(n1746), .B0(n5355), .B1(n7389), .C0(n1762), 
        .Y(n3622) );
  NAND2X1 U6828 ( .A(N7688), .B(n7218), .Y(n1762) );
  OAI221X1 U6829 ( .A0(n7604), .A1(n1746), .B0(n5355), .B1(n7390), .C0(n1760), 
        .Y(n3621) );
  NAND2X1 U6830 ( .A(N7689), .B(n7218), .Y(n1760) );
  OAI221X1 U6831 ( .A0(n7605), .A1(n1746), .B0(n5355), .B1(n7391), .C0(n1758), 
        .Y(n3620) );
  NAND2X1 U6832 ( .A(N7690), .B(n7218), .Y(n1758) );
  NOR2X1 U6833 ( .A(n1910), .B(n2153), .Y(n5013) );
  OAI221X1 U6834 ( .A0(n2154), .A1(n7206), .B0(n6239), .B1(n6776), .C0(n6238), 
        .Y(n6286) );
  AOI211X1 U6835 ( .A0(n7032), .A1(n7326), .B0(n7012), .C0(n5013), .Y(n2154)
         );
  AOI31X1 U6836 ( .A0(n7030), .A1(n6237), .A2(n1910), .B0(n5350), .Y(n6238) );
  INVX2 U6837 ( .A(n2153), .Y(n6237) );
  OR4X2 U6838 ( .A(n818), .B(n7247), .C(n819), .D(n837), .Y(n878) );
  INVX2 U6839 ( .A(N7477), .Y(n5075) );
  NAND3X1 U6840 ( .A(n1909), .B(n7033), .C(n6092), .Y(n6138) );
  AOI31X1 U6841 ( .A0(n7328), .A1(n1910), .A2(n7024), .B0(n1911), .Y(n1909) );
  AOI32X1 U6842 ( .A0(n6498), .A1(n2106), .A2(n7324), .B0(n1907), .B1(n7034), 
        .Y(n6092) );
  INVX2 U6843 ( .A(n6792), .Y(n7024) );
  OAI211X1 U6844 ( .A0(n1910), .A1(n6391), .B0(n4850), .C0(n7033), .Y(n6441)
         );
  INVX2 U6845 ( .A(n6032), .Y(N7433) );
  OAI221X1 U6846 ( .A0(n7609), .A1(n1831), .B0(n7197), .B1(n7396), .C0(n1845), 
        .Y(n3676) );
  NAND2X1 U6847 ( .A(N7648), .B(n7195), .Y(n1845) );
  OAI221X1 U6848 ( .A0(n7610), .A1(n1831), .B0(n7197), .B1(n7397), .C0(n1843), 
        .Y(n3675) );
  NAND2X1 U6849 ( .A(N7649), .B(n7195), .Y(n1843) );
  OAI221X1 U6850 ( .A0(n7611), .A1(n1831), .B0(n7197), .B1(n7394), .C0(n1841), 
        .Y(n3674) );
  NAND2X1 U6851 ( .A(N7650), .B(n7195), .Y(n1841) );
  OAI222X1 U6852 ( .A0(n5024), .A1(n1435), .B0(n7558), .B1(n1436), .C0(n4850), 
        .C1(n7368), .Y(n3287) );
  OAI222X1 U6853 ( .A0(n7552), .A1(n1435), .B0(n7556), .B1(n1436), .C0(n4850), 
        .C1(n7364), .Y(n3289) );
  OAI222X1 U6854 ( .A0(n7553), .A1(n1435), .B0(n7557), .B1(n1436), .C0(n4850), 
        .C1(n7369), .Y(n3288) );
  OAI222X1 U6855 ( .A0(n5365), .A1(n1435), .B0(N7907), .B1(n1436), .C0(n4850), 
        .C1(n7365), .Y(n3292) );
  OAI221X1 U6856 ( .A0(n7613), .A1(n1831), .B0(n7197), .B1(n7398), .C0(n1834), 
        .Y(n3672) );
  NAND2X1 U6857 ( .A(N7652), .B(n7195), .Y(n1834) );
  OAI221X1 U6858 ( .A0(n7612), .A1(n1831), .B0(n7197), .B1(n7399), .C0(n1838), 
        .Y(n3673) );
  NAND2X1 U6859 ( .A(N7651), .B(n7195), .Y(n1838) );
  OAI221X1 U6860 ( .A0(N7475), .A1(n2156), .B0(n5351), .B1(n7431), .C0(n2172), 
        .Y(n3897) );
  NAND2X1 U6861 ( .A(N7475), .B(n7209), .Y(n2172) );
  OAI221X1 U6862 ( .A0(n7630), .A1(n2156), .B0(n5351), .B1(n7432), .C0(n2170), 
        .Y(n3896) );
  NAND2X1 U6863 ( .A(N7476), .B(n7209), .Y(n2170) );
  OAI221X1 U6864 ( .A0(n7631), .A1(n2156), .B0(n5351), .B1(n7433), .C0(n2168), 
        .Y(n3895) );
  NAND2X1 U6865 ( .A(N7477), .B(n7209), .Y(n2168) );
  OAI222X1 U6866 ( .A0(n7543), .A1(n1381), .B0(n7546), .B1(n1383), .C0(n4847), 
        .C1(n7343), .Y(n3235) );
  INVX2 U6867 ( .A(n6040), .Y(N7434) );
  OR2X1 U6868 ( .A(n5374), .B(n7230), .Y(n6792) );
  OAI211X1 U6869 ( .A0(n6721), .A1(n6792), .B0(n6720), .C0(n7033), .Y(n6771)
         );
  INVX2 U6870 ( .A(N7567), .Y(n5165) );
  INVX2 U6871 ( .A(N7947), .Y(n7545) );
  OAI221X1 U6872 ( .A0(n4934), .A1(n1831), .B0(n7197), .B1(n7395), .C0(n1847), 
        .Y(n3677) );
  NAND2X1 U6873 ( .A(n4934), .B(n7195), .Y(n1847) );
  OAI2BB1X1 U6874 ( .A0N(n7028), .A1N(n5376), .B0(n5903), .Y(n6030) );
  OAI2BB1X1 U6875 ( .A0N(n7230), .A1N(n7206), .B0(n5006), .Y(n5903) );
  OAI221X1 U6876 ( .A0(N7565), .A1(n1994), .B0(n5353), .B1(n7411), .C0(n2011), 
        .Y(n3787) );
  NAND2X1 U6877 ( .A(N7565), .B(n7214), .Y(n2011) );
  OAI211X1 U6878 ( .A0(n6609), .A1(n6792), .B0(n6608), .C0(n7033), .Y(n6661)
         );
  AOI2BB2X1 U6879 ( .B0(n7015), .B1(n7038), .A0N(n7035), .A1N(n1585), .Y(n6609) );
  OAI221X1 U6880 ( .A0(n7621), .A1(n1994), .B0(n5353), .B1(n7410), .C0(n2002), 
        .Y(n3784) );
  NAND2X1 U6881 ( .A(N7568), .B(n7214), .Y(n2002) );
  OAI221X1 U6882 ( .A0(n7623), .A1(n1994), .B0(n5353), .B1(n7414), .C0(n1997), 
        .Y(n3782) );
  NAND2X1 U6883 ( .A(N7570), .B(n7214), .Y(n1997) );
  OAI221X1 U6884 ( .A0(n7622), .A1(n1994), .B0(n5353), .B1(n7415), .C0(n2000), 
        .Y(n3783) );
  NAND2X1 U6885 ( .A(N7569), .B(n7214), .Y(n2000) );
  NOR4BX1 U6886 ( .AN(n2809), .B(n5006), .C(n7020), .D(n7321), .Y(n2776) );
  AOI221XL U6887 ( .A0(n2710), .A1(n7021), .B0(n2810), .B1(n7328), .C0(n2731), 
        .Y(n2809) );
  NOR2X1 U6888 ( .A(n5376), .B(n2708), .Y(n2810) );
  OR2X1 U6889 ( .A(n2153), .B(n2804), .Y(n6774) );
  INVX2 U6890 ( .A(N7839), .Y(n7572) );
  OAI31X1 U6891 ( .A0(n2697), .A1(n2696), .A2(n6776), .B0(n2783), .Y(n2748) );
  OAI221X1 U6892 ( .A0(N7521), .A1(n2075), .B0(n7213), .B1(n7422), .C0(n2090), 
        .Y(n3842) );
  NAND2X1 U6893 ( .A(N7521), .B(n7211), .Y(n2090) );
  OAI221X1 U6894 ( .A0(N7606), .A1(n1913), .B0(n5354), .B1(n7403), .C0(n1929), 
        .Y(n3732) );
  NAND2X1 U6895 ( .A(N7606), .B(n7216), .Y(n1929) );
  OAI222X1 U6896 ( .A0(n5364), .A1(n1536), .B0(N7835), .B1(n1538), .C0(n5358), 
        .C1(n7347), .Y(n3402) );
  OAI222X1 U6897 ( .A0(n7542), .A1(n1381), .B0(n4901), .B1(n1383), .C0(n4847), 
        .C1(n7342), .Y(n3236) );
  INVX2 U6898 ( .A(N7944), .Y(n7542) );
  OAI222X1 U6899 ( .A0(n7571), .A1(n1536), .B0(n7577), .B1(n1538), .C0(n5358), 
        .C1(n7350), .Y(n3397) );
  OAI222X1 U6900 ( .A0(n7572), .A1(n1536), .B0(n7576), .B1(n1538), .C0(n5358), 
        .C1(n7351), .Y(n3398) );
  OAI222X1 U6901 ( .A0(n7570), .A1(n1536), .B0(n7575), .B1(n1538), .C0(n5358), 
        .C1(n7346), .Y(n3399) );
  OAI222X1 U6902 ( .A0(n7569), .A1(n1536), .B0(n7574), .B1(n1538), .C0(n5358), 
        .C1(n7349), .Y(n3400) );
  OAI222X1 U6903 ( .A0(n7568), .A1(n1536), .B0(n7573), .B1(n1538), .C0(n5358), 
        .C1(n7348), .Y(n3401) );
  INVX2 U6904 ( .A(N7836), .Y(n7568) );
  OAI222X1 U6905 ( .A0(n7597), .A1(n1691), .B0(n7601), .B1(n1693), .C0(n5356), 
        .C1(n7382), .Y(n3565) );
  OAI222X1 U6906 ( .A0(n7596), .A1(n1691), .B0(n7600), .B1(n1693), .C0(n5356), 
        .C1(n7381), .Y(n3566) );
  INVX2 U6907 ( .A(N7728), .Y(n7596) );
  OAI222X1 U6908 ( .A0(n5018), .A1(n1642), .B0(n7595), .B1(n1643), .C0(n5357), 
        .C1(n7362), .Y(n3507) );
  OAI222X1 U6909 ( .A0(n7590), .A1(n1642), .B0(n7594), .B1(n1643), .C0(n5357), 
        .C1(n7363), .Y(n3508) );
  OAI222X1 U6910 ( .A0(n7589), .A1(n1642), .B0(n7593), .B1(n1643), .C0(n5357), 
        .C1(n7358), .Y(n3509) );
  OAI222X1 U6911 ( .A0(n7588), .A1(n1642), .B0(n7592), .B1(n1643), .C0(n5357), 
        .C1(n7361), .Y(n3510) );
  OAI222X1 U6912 ( .A0(n7587), .A1(n1642), .B0(n7591), .B1(n1643), .C0(n5357), 
        .C1(n7360), .Y(n3511) );
  INVX2 U6913 ( .A(N7764), .Y(n7587) );
  OAI222X1 U6914 ( .A0(n7579), .A1(n1587), .B0(n7583), .B1(n1589), .C0(n4851), 
        .C1(n7355), .Y(n3455) );
  OAI222X1 U6915 ( .A0(n7578), .A1(n1587), .B0(n7582), .B1(n1589), .C0(n4851), 
        .C1(n7354), .Y(n3456) );
  INVX2 U6916 ( .A(N7800), .Y(n7578) );
  OAI222X1 U6917 ( .A0(n7560), .A1(n1486), .B0(n7564), .B1(n1488), .C0(n5359), 
        .C1(n7373), .Y(n3345) );
  OAI222X1 U6918 ( .A0(n7559), .A1(n1486), .B0(n7563), .B1(n1488), .C0(n5359), 
        .C1(n7372), .Y(n3346) );
  INVX2 U6919 ( .A(N7872), .Y(n7559) );
  OAI222X1 U6920 ( .A0(n5028), .A1(n1587), .B0(n7586), .B1(n1589), .C0(n4851), 
        .C1(n7356), .Y(n3452) );
  OAI222X1 U6921 ( .A0(n7581), .A1(n1587), .B0(n7585), .B1(n1589), .C0(n4851), 
        .C1(n7357), .Y(n3453) );
  OAI222X1 U6922 ( .A0(n7580), .A1(n1587), .B0(n7584), .B1(n1589), .C0(n4851), 
        .C1(n7352), .Y(n3454) );
  OAI221X1 U6923 ( .A0(n7625), .A1(n2075), .B0(n7213), .B1(n7423), .C0(n2088), 
        .Y(n3841) );
  NAND2X1 U6924 ( .A(N7522), .B(n7211), .Y(n2088) );
  OAI221X1 U6925 ( .A0(n7626), .A1(n2075), .B0(n7213), .B1(n7424), .C0(n2086), 
        .Y(n3840) );
  NAND2X1 U6926 ( .A(N7523), .B(n7211), .Y(n2086) );
  OAI221X1 U6927 ( .A0(n7627), .A1(n2075), .B0(n7213), .B1(n7421), .C0(n2084), 
        .Y(n3839) );
  NAND2X1 U6928 ( .A(N7524), .B(n7211), .Y(n2084) );
  OAI221X1 U6929 ( .A0(n7629), .A1(n2075), .B0(n7213), .B1(n7425), .C0(n2078), 
        .Y(n3837) );
  NAND2X1 U6930 ( .A(N7526), .B(n7211), .Y(n2078) );
  OAI221X1 U6931 ( .A0(n7628), .A1(n2075), .B0(n7213), .B1(n7426), .C0(n2082), 
        .Y(n3838) );
  NAND2X1 U6932 ( .A(N7525), .B(n7211), .Y(n2082) );
  NOR2X1 U6933 ( .A(n5573), .B(n5572), .Y(n2733) );
  OR2X1 U6934 ( .A(n6780), .B(n6789), .Y(n835) );
  OAI222X1 U6935 ( .A0(n5016), .A1(n1327), .B0(n7541), .B1(n1328), .C0(n5360), 
        .C1(n7338), .Y(n3177) );
  OAI222X1 U6936 ( .A0(n7535), .A1(n1327), .B0(n7539), .B1(n1328), .C0(n5360), 
        .C1(n7334), .Y(n3179) );
  OAI222X1 U6937 ( .A0(n7534), .A1(n1327), .B0(n7538), .B1(n1328), .C0(n5360), 
        .C1(n7337), .Y(n3180) );
  OAI222X1 U6938 ( .A0(n7533), .A1(n1327), .B0(n7537), .B1(n1328), .C0(n5360), 
        .C1(n7336), .Y(n3181) );
  INVX2 U6939 ( .A(N7980), .Y(n7533) );
  OAI222X1 U6940 ( .A0(n7536), .A1(n1327), .B0(n7540), .B1(n1328), .C0(n5360), 
        .C1(n7339), .Y(n3178) );
  NOR2X1 U6941 ( .A(n7206), .B(n2789), .Y(n2772) );
  AOI221XL U6942 ( .A0(n5374), .A1(n2701), .B0(n7329), .B1(n7324), .C0(n7327), 
        .Y(n2789) );
  OAI2BB1X1 U6943 ( .A0N(n2788), .A1N(n1910), .B0(n2772), .Y(n2765) );
  INVX2 U6944 ( .A(N7911), .Y(n7553) );
  OAI221X1 U6945 ( .A0(n7614), .A1(n1913), .B0(n5354), .B1(n7404), .C0(n1927), 
        .Y(n3731) );
  NAND2X1 U6946 ( .A(N7607), .B(n7216), .Y(n1927) );
  OAI221X1 U6947 ( .A0(n7615), .A1(n1913), .B0(n5354), .B1(n7405), .C0(n1925), 
        .Y(n3730) );
  NAND2X1 U6948 ( .A(N7608), .B(n7216), .Y(n1925) );
  INVX2 U6949 ( .A(N7731), .Y(n7599) );
  INVX2 U6950 ( .A(N7803), .Y(n7581) );
  INVX2 U6951 ( .A(n5572), .Y(n5571) );
  NAND3X1 U6952 ( .A(n7033), .B(n2388), .C(n2389), .Y(n2366) );
  NAND4X1 U6953 ( .A(n2468), .B(n2469), .C(n2470), .D(n2471), .Y(n2394) );
  AOI222XL U6954 ( .A0(n2485), .A1(n7011), .B0(n2487), .B1(n2488), .C0(n2489), 
        .C1(n2490), .Y(n2470) );
  AOI221XL U6955 ( .A0(n2472), .A1(n2473), .B0(n2474), .B1(n2475), .C0(n2476), 
        .Y(n2471) );
  AOI222XL U6956 ( .A0(n2508), .A1(n2509), .B0(n2510), .B1(n2511), .C0(n2512), 
        .C1(n2513), .Y(n2468) );
  OAI2BB2X1 U6957 ( .B0(n7292), .B1(n2366), .A0N(N8519), .A1N(n7204), .Y(n4008) );
  OAI2BB2X1 U6958 ( .B0(n7270), .B1(n2366), .A0N(N8518), .A1N(n7204), .Y(n4027) );
  NAND2BX1 U6959 ( .AN(n2775), .B(n2776), .Y(n2758) );
  INVX2 U6960 ( .A(n875), .Y(n7282) );
  NOR2X1 U6961 ( .A(n2397), .B(n831), .Y(n1350) );
  OAI2BB2X1 U6962 ( .B0(n4849), .B1(n2366), .A0N(N8520), .A1N(n7204), .Y(n4007) );
  NAND4X1 U6963 ( .A(n2405), .B(n2406), .C(n2407), .D(n2408), .Y(n2392) );
  AOI32X1 U6964 ( .A0(n2099), .A1(n7500), .A2(n2100), .B0(n2409), .B1(n2410), 
        .Y(n2408) );
  AOI33X1 U6965 ( .A0(n1856), .A1(n7523), .A2(n1857), .B0(n7263), .B1(n7497), 
        .B2(n1772), .Y(n2406) );
  AOI33X1 U6966 ( .A0(n7274), .A1(n7418), .A2(n2021), .B0(n7276), .B1(n7513), 
        .B2(n1939), .Y(n2407) );
  AOI33X1 U6967 ( .A0(n7273), .A1(n7385), .A2(n1712), .B0(n7278), .B1(n7510), 
        .B2(n1660), .Y(n2405) );
  INVX2 U6968 ( .A(n1713), .Y(n7273) );
  OAI22X1 U6969 ( .A0(n5361), .A1(n7626), .B0(n188), .B1(n7627), .Y(n768) );
  NOR2X1 U6970 ( .A(n5415), .B(n745), .Y(n2265) );
  OAI22X1 U6971 ( .A0(N11045), .A1(n93), .B0(n94), .B1(n7298), .Y(
        next_state[1]) );
  OAI222X1 U6972 ( .A0(n745), .A1(n188), .B0(n193), .B1(n884), .C0(n5362), 
        .C1(n867), .Y(n819) );
  INVX2 U6973 ( .A(n2388), .Y(n7204) );
  NAND4X1 U6974 ( .A(n5364), .B(n7265), .C(n2401), .D(n7573), .Y(n2478) );
  OAI22X1 U6975 ( .A0(n4851), .A1(n7354), .B0(n1609), .B1(n4898), .Y(n3465) );
  NAND2BX1 U6976 ( .AN(n2459), .B(n2389), .Y(n2458) );
  NAND4BX1 U6977 ( .AN(n2462), .B(n2463), .C(n2464), .D(n2465), .Y(n2459) );
  AOI33X1 U6978 ( .A0(n7265), .A1(n7494), .A2(n1556), .B0(n7272), .B1(n7376), 
        .B2(n1507), .Y(n2463) );
  AOI33X1 U6979 ( .A0(n7279), .A1(n7510), .A2(n1660), .B0(n199), .B1(n7520), 
        .B2(n1607), .Y(n2464) );
  NAND4BX1 U6980 ( .AN(n2527), .B(n2528), .C(n2529), .D(n2530), .Y(n2462) );
  NOR2X1 U6981 ( .A(n7532), .B(n2458), .Y(N8757) );
  NOR2X1 U6982 ( .A(n7531), .B(n2458), .Y(N8756) );
  NOR2X1 U6983 ( .A(n7530), .B(n2458), .Y(N8755) );
  NOR2X1 U6984 ( .A(n7529), .B(n2458), .Y(N8754) );
  NOR2X1 U6985 ( .A(n7259), .B(n2458), .Y(N8753) );
  AOI33X1 U6986 ( .A0(n7271), .A1(n7376), .A2(n1507), .B0(n7289), .B1(n7516), 
        .B2(n7518), .Y(n2399) );
  INVX2 U6987 ( .A(n1402), .Y(n7289) );
  INVX2 U6988 ( .A(N7431), .Y(n5344) );
  NAND2X1 U6989 ( .A(n2415), .B(n7275), .Y(n2022) );
  NAND2X1 U6990 ( .A(n2418), .B(n7279), .Y(n1661) );
  OAI22X1 U6991 ( .A0(n5355), .A1(n7391), .B0(n1774), .B1(n4948), .Y(n3629) );
  OAI22X1 U6992 ( .A0(n5355), .A1(n7390), .B0(n1774), .B1(n4896), .Y(n3630) );
  INVX2 U6993 ( .A(n1773), .Y(n7263) );
  NOR2X1 U6994 ( .A(n2401), .B(n182), .Y(n1555) );
  AOI33X1 U6995 ( .A0(n7288), .A1(n7520), .A2(n1607), .B0(n1555), .B1(n7494), 
        .B2(n1556), .Y(n2400) );
  NAND3X1 U6996 ( .A(n7622), .B(n7623), .C(n7621), .Y(n913) );
  OAI22X1 U6997 ( .A0(n5356), .A1(n7381), .B0(n1714), .B1(n4892), .Y(n3575) );
  OAI22X1 U6998 ( .A0(n5359), .A1(n7372), .B0(n1509), .B1(n4899), .Y(n3355) );
  OAI22X1 U6999 ( .A0(n4850), .A1(n7366), .B0(n1457), .B1(n4895), .Y(n3300) );
  OAI22X1 U7000 ( .A0(n5357), .A1(n7360), .B0(n1662), .B1(n4894), .Y(n3520) );
  OAI22X1 U7001 ( .A0(n4847), .A1(n7342), .B0(n1404), .B1(n4893), .Y(n3245) );
  OAI22X1 U7002 ( .A0(n5360), .A1(n7336), .B0(n1351), .B1(n4900), .Y(n3190) );
  NOR4X1 U7003 ( .A(n928), .B(n2412), .C(n831), .D(n4952), .Y(n2409) );
  NAND2X1 U7004 ( .A(n929), .B(n2397), .Y(n2412) );
  NAND2X1 U7005 ( .A(n2398), .B(n7281), .Y(n1456) );
  OAI22X1 U7006 ( .A0(n5358), .A1(n7348), .B0(n1558), .B1(n4897), .Y(n3410) );
  INVX2 U7007 ( .A(n5569), .Y(n5568) );
  OAI22X1 U7008 ( .A0(n7197), .A1(n7397), .B0(n1859), .B1(n7401), .Y(n3684) );
  OAI22X1 U7009 ( .A0(n7197), .A1(n7396), .B0(n1859), .B1(n7400), .Y(n3685) );
  NAND2X1 U7010 ( .A(n2414), .B(n7277), .Y(n1940) );
  OAI22X1 U7011 ( .A0(n5351), .A1(n7433), .B0(n2276), .B1(n7437), .Y(n3983) );
  OAI22X1 U7012 ( .A0(n5351), .A1(n7432), .B0(n2276), .B1(n7436), .Y(n3982) );
  AND2X1 U7013 ( .A(n2459), .B(n2389), .Y(N8752) );
  OAI211X1 U7014 ( .A0(n2750), .A1(n7234), .B0(n2762), .C0(n2763), .Y(n2761)
         );
  OAI22X1 U7015 ( .A0(n2102), .A1(n7428), .B0(n7213), .B1(n7423), .Y(n3850) );
  OAI22X1 U7016 ( .A0(n188), .A1(n7556), .B0(n190), .B1(n7558), .Y(n187) );
  NAND2BX1 U7017 ( .AN(n2402), .B(n199), .Y(n1608) );
  OAI22X1 U7018 ( .A0(n5353), .A1(n7412), .B0(n2023), .B1(n7416), .Y(n3795) );
  OAI22X1 U7019 ( .A0(n5353), .A1(n7413), .B0(n2023), .B1(n7417), .Y(n3794) );
  INVX2 U7020 ( .A(N7419), .Y(n7047) );
  OAI22X1 U7021 ( .A0(n5354), .A1(n7404), .B0(n1941), .B1(n7408), .Y(n3740) );
  NAND2X1 U7022 ( .A(n2404), .B(n7272), .Y(n1508) );
  NOR2X1 U7023 ( .A(n2413), .B(n761), .Y(n2099) );
  OAI22X1 U7024 ( .A0(n4850), .A1(n7367), .B0(n1457), .B1(n4947), .Y(n3299) );
  OAI22X1 U7025 ( .A0(n2102), .A1(n7429), .B0(n7213), .B1(n7424), .Y(n3849) );
  NOR2X1 U7026 ( .A(n2417), .B(n882), .Y(n1856) );
  OAI22X1 U7027 ( .A0(n4847), .A1(n7343), .B0(n1404), .B1(n4945), .Y(n3244) );
  OAI22X1 U7028 ( .A0(n5354), .A1(n7405), .B0(n1941), .B1(n7409), .Y(n3739) );
  OAI22X1 U7029 ( .A0(n868), .A1(n882), .B0(n883), .B1(n884), .Y(n880) );
  NOR2X1 U7030 ( .A(n7260), .B(n836), .Y(n883) );
  OAI22X1 U7031 ( .A0(n5358), .A1(n7349), .B0(n1558), .B1(n4949), .Y(n3409) );
  OAI22X1 U7032 ( .A0(n5356), .A1(n7382), .B0(n1714), .B1(n4944), .Y(n3574) );
  OAI22X1 U7033 ( .A0(n5357), .A1(n7361), .B0(n1662), .B1(n4946), .Y(n3519) );
  OR2X1 U7034 ( .A(n7039), .B(n6390), .Y(n6793) );
  OAI22X1 U7035 ( .A0(n5359), .A1(n7373), .B0(n1509), .B1(n4951), .Y(n3354) );
  OAI22X1 U7036 ( .A0(n4851), .A1(n7355), .B0(n1609), .B1(n4950), .Y(n3464) );
  OAI22X1 U7037 ( .A0(n5360), .A1(n7337), .B0(n1351), .B1(n4953), .Y(n3189) );
  AOI33X1 U7038 ( .A0(n1712), .A1(n7385), .A2(n5015), .B0(n1772), .B1(n7497), 
        .B2(n7264), .Y(n2530) );
  NOR2X1 U7039 ( .A(n1314), .B(n5464), .Y(n2436) );
  AND3X2 U7040 ( .A(n2436), .B(n7301), .C(n5572), .Y(n2454) );
  AOI33X1 U7041 ( .A0(n2021), .A1(n7418), .A2(n7275), .B0(n2100), .B1(n7500), 
        .B2(n7261), .Y(n2528) );
  NAND3X1 U7042 ( .A(n7540), .B(n7541), .C(n7539), .Y(n832) );
  NOR2X1 U7043 ( .A(n1314), .B(n5442), .Y(n2433) );
  AND3X2 U7044 ( .A(n2433), .B(n5570), .C(n2431), .Y(n2435) );
  INVX2 U7045 ( .A(n96), .Y(n5900) );
  NAND2X1 U7046 ( .A(n7261), .B(n876), .Y(n873) );
  AOI33X1 U7047 ( .A0(n1857), .A1(n7523), .A2(n7286), .B0(n1939), .B1(n7513), 
        .B2(n7277), .Y(n2529) );
  NAND2X1 U7048 ( .A(n2420), .B(n7285), .Y(n2272) );
  NAND2X1 U7049 ( .A(n7309), .B(n5573), .Y(n2430) );
  AOI32X1 U7050 ( .A0(n5571), .A1(n5570), .A2(n2430), .B0(n5014), .B1(N5061), 
        .Y(n2432) );
  AND2X1 U7051 ( .A(n7308), .B(n5572), .Y(n5014) );
  INVX2 U7052 ( .A(n6789), .Y(n7011) );
  AOI33X1 U7053 ( .A0(n2431), .A1(n2433), .A2(n2447), .B0(n2436), .B1(n2445), 
        .B2(n2448), .Y(WEN23) );
  NOR2X1 U7054 ( .A(n2442), .B(n5570), .Y(n2447) );
  OAI21X1 U7055 ( .A0(n7516), .A1(n1403), .B0(n1395), .Y(n1398) );
  NAND4X1 U7056 ( .A(n7303), .B(n7302), .C(n7304), .D(n7305), .Y(n2439) );
  INVX2 U7057 ( .A(n2493), .Y(n6781) );
  OAI21X1 U7058 ( .A0(n7503), .A1(n1348), .B0(n1342), .Y(n1345) );
  NAND2X1 U7059 ( .A(n2397), .B(n7537), .Y(n2522) );
  OAI21X1 U7060 ( .A0(n7526), .A1(n2273), .B0(n2267), .Y(n2270) );
  NAND2X1 U7061 ( .A(n5014), .B(n5570), .Y(n104) );
  AOI22X1 U7062 ( .A0(n2436), .A1(n7299), .B0(n2433), .B1(n2438), .Y(WEN33) );
  INVX2 U7063 ( .A(n2444), .Y(n7299) );
  OAI33X1 U7064 ( .A0(n5569), .A1(n2439), .A2(n104), .B0(n2440), .B1(n7308), 
        .B2(n2442), .Y(n2438) );
  AOI32X1 U7065 ( .A0(n2445), .A1(n2446), .A2(N5059), .B0(n7301), .B1(n5014), 
        .Y(n2444) );
  NAND2X1 U7066 ( .A(n5457), .B(n5567), .Y(n119) );
  INVX2 U7067 ( .A(n1403), .Y(n7518) );
  INVX2 U7068 ( .A(length9[4]), .Y(n7357) );
  NOR2X1 U7069 ( .A(n7509), .B(n7508), .Y(n1455) );
  NOR2X1 U7070 ( .A(n7515), .B(n7514), .Y(n1939) );
  NOR2X1 U7071 ( .A(n5572), .B(n2439), .Y(n2445) );
  NAND3X1 U7072 ( .A(n7557), .B(n7558), .C(n7556), .Y(n809) );
  NOR2X1 U7073 ( .A(n7499), .B(n7498), .Y(n1772) );
  NOR2X1 U7074 ( .A(n7502), .B(n7501), .Y(n2100) );
  NOR2X1 U7075 ( .A(n7512), .B(n7511), .Y(n1660) );
  NOR3X1 U7076 ( .A(n2439), .B(n5415), .C(n1314), .Y(n2449) );
  NOR2X1 U7077 ( .A(n7496), .B(n7495), .Y(n1556) );
  NOR2X1 U7078 ( .A(n7420), .B(n7419), .Y(n2021) );
  NOR2X1 U7079 ( .A(n7525), .B(n7524), .Y(n1857) );
  NOR2X1 U7080 ( .A(n7387), .B(n7386), .Y(n1712) );
  NOR2X1 U7081 ( .A(n7522), .B(n7521), .Y(n1607) );
  NOR2X1 U7082 ( .A(n7378), .B(n7377), .Y(n1507) );
  XOR2X1 U7083 ( .A(n5573), .B(n7309), .Y(n2448) );
  NAND2X1 U7084 ( .A(n7301), .B(n5569), .Y(n2442) );
  INVX2 U7085 ( .A(n111), .Y(n5466) );
  NOR2X1 U7086 ( .A(n5374), .B(n5376), .Y(n1829) );
  BUFX2 U7087 ( .A(n1340), .Y(n5352) );
  NOR3BX1 U7088 ( .AN(n929), .B(n96), .C(n928), .Y(n1340) );
  INVX2 U7089 ( .A(length7[4]), .Y(n7384) );
  INVX2 U7090 ( .A(length10[4]), .Y(n7351) );
  INVX2 U7091 ( .A(length13[4]), .Y(n7345) );
  INVX2 U7092 ( .A(length14[4]), .Y(n7339) );
  INVX2 U7093 ( .A(length11[4]), .Y(n7375) );
  INVX2 U7094 ( .A(length12[4]), .Y(n7369) );
  INVX2 U7095 ( .A(length8[4]), .Y(n7363) );
  INVX2 U7096 ( .A(length9[5]), .Y(n7356) );
  NAND2X1 U7097 ( .A(n5466), .B(n5567), .Y(n118) );
  INVX2 U7098 ( .A(n102), .Y(n7297) );
  INVX2 U7099 ( .A(length5[4]), .Y(n7399) );
  INVX2 U7100 ( .A(length1[4]), .Y(n7435) );
  INVX2 U7101 ( .A(length2[4]), .Y(n7426) );
  INVX2 U7102 ( .A(length3[4]), .Y(n7415) );
  INVX2 U7103 ( .A(length4[4]), .Y(n7407) );
  INVX2 U7104 ( .A(length6[4]), .Y(n7393) );
  INVX2 U7105 ( .A(n5378), .Y(n7312) );
  INVX2 U7106 ( .A(n7232), .Y(n5436) );
  INVX2 U7107 ( .A(length10[5]), .Y(n7350) );
  INVX2 U7108 ( .A(length11[5]), .Y(n7374) );
  INVX2 U7109 ( .A(length12[5]), .Y(n7368) );
  INVX2 U7110 ( .A(length8[5]), .Y(n7362) );
  INVX2 U7111 ( .A(length13[5]), .Y(n7344) );
  INVX2 U7112 ( .A(length14[5]), .Y(n7338) );
  INVX2 U7113 ( .A(length7[5]), .Y(n7383) );
  NOR2X1 U7114 ( .A(n5570), .B(n5572), .Y(n1270) );
  INVX2 U7115 ( .A(length1[5]), .Y(n7434) );
  INVX2 U7116 ( .A(length2[5]), .Y(n7425) );
  INVX2 U7117 ( .A(length3[5]), .Y(n7414) );
  INVX2 U7118 ( .A(length4[5]), .Y(n7406) );
  INVX2 U7119 ( .A(length5[5]), .Y(n7398) );
  INVX2 U7120 ( .A(length6[5]), .Y(n7392) );
  OAI2BB1X1 U7121 ( .A0N(N5804), .A1N(n4991), .B0(n6093), .Y(n3726) );
  OAI2BB1X1 U7122 ( .A0N(N5541), .A1N(n5002), .B0(n6240), .Y(n3891) );
  OR2X1 U7123 ( .A(n6606), .B(n6605), .Y(n6607) );
  OR2X1 U7124 ( .A(n6717), .B(n6716), .Y(n6718) );
  OAI2BB1X1 U7125 ( .A0N(N5539), .A1N(n5002), .B0(n6242), .Y(n3853) );
  OAI2BB1X1 U7126 ( .A0N(N5802), .A1N(n4991), .B0(n6095), .Y(n3688) );
  OR2X1 U7127 ( .A(n6388), .B(n6387), .Y(n6389) );
  OAI2BB1XL U7128 ( .A0N(N6292), .A1N(n4996), .B0(n6663), .Y(n3506) );
  OR2X1 U7129 ( .A(n6662), .B(n6661), .Y(n6663) );
  OAI2BB1X1 U7130 ( .A0N(N5722), .A1N(n4998), .B0(n6190), .Y(n3836) );
  OR2X1 U7131 ( .A(n6772), .B(n6771), .Y(n6773) );
  OAI2BB1X1 U7132 ( .A0N(N5763), .A1N(n4989), .B0(n6141), .Y(n3781) );
  OR2X1 U7133 ( .A(n6496), .B(n6495), .Y(n6497) );
  OAI2BB1X1 U7134 ( .A0N(N5500), .A1N(n5003), .B0(n6291), .Y(n3937) );
  OR2X1 U7135 ( .A(n6442), .B(n6441), .Y(n6443) );
  OAI2BB1X1 U7136 ( .A0N(N5459), .A1N(n5005), .B0(n5904), .Y(n3977) );
  OR2X1 U7137 ( .A(n6550), .B(n6549), .Y(n6551) );
  OAI2BB1X1 U7138 ( .A0N(N5803), .A1N(n4991), .B0(n6094), .Y(n3687) );
  OAI2BB1X1 U7139 ( .A0N(N5540), .A1N(n5002), .B0(n6241), .Y(n3852) );
  OAI2BB1X1 U7140 ( .A0N(N5761), .A1N(n4989), .B0(n6143), .Y(n3743) );
  AND3X2 U7141 ( .A(n7008), .B(n5400), .C(n7006), .Y(n7009) );
  INVX2 U7142 ( .A(n7002), .Y(n7008) );
  AOI222XL U7143 ( .A0(reg_length0[4]), .A1(n7018), .B0(reg_length0[0]), .B1(
        n7012), .C0(reg_length0[3]), .C1(n5013), .Y(n6990) );
  OR2X1 U7144 ( .A(n6553), .B(n6605), .Y(n6554) );
  OAI2BB1X1 U7145 ( .A0N(N5457), .A1N(n5005), .B0(n5906), .Y(n3939) );
  OAI2BB1X1 U7146 ( .A0N(N5721), .A1N(n4998), .B0(n6191), .Y(n3797) );
  OAI2BB1X1 U7147 ( .A0N(N5843), .A1N(n4990), .B0(n6047), .Y(n3633) );
  OAI2BB1X1 U7148 ( .A0N(N5538), .A1N(n5002), .B0(n6243), .Y(n3854) );
  OAI2BB1X1 U7149 ( .A0N(N5801), .A1N(n4991), .B0(n6096), .Y(n3689) );
  OAI2BB1X1 U7150 ( .A0N(N5458), .A1N(n5005), .B0(n5905), .Y(n3938) );
  OAI2BB1X1 U7151 ( .A0N(N5498), .A1N(n5003), .B0(n6293), .Y(n3899) );
  OAI2BB1X1 U7152 ( .A0N(N5499), .A1N(n5003), .B0(n6292), .Y(n3898) );
  OAI2BB1X1 U7153 ( .A0N(N5720), .A1N(n4998), .B0(n6192), .Y(n3798) );
  OAI2BB1X1 U7154 ( .A0N(N5452), .A1N(n5005), .B0(n5911), .Y(n3944) );
  OAI2BB1X1 U7155 ( .A0N(N5451), .A1N(n5005), .B0(n5912), .Y(n3945) );
  OAI2BB1X1 U7156 ( .A0N(N5453), .A1N(n5005), .B0(n5910), .Y(n3943) );
  OAI2BB1X1 U7157 ( .A0N(N5454), .A1N(n5005), .B0(n5909), .Y(n3942) );
  OAI2BB1X1 U7158 ( .A0N(N5456), .A1N(n5005), .B0(n5907), .Y(n3940) );
  OAI2BB1X1 U7159 ( .A0N(N5455), .A1N(n5005), .B0(n5908), .Y(n3941) );
  OAI2BB1X1 U7160 ( .A0N(N5840), .A1N(n4990), .B0(n6050), .Y(n3636) );
  OAI2BB1X1 U7161 ( .A0N(N5760), .A1N(n4989), .B0(n6144), .Y(n3744) );
  OAI2BB1X1 U7162 ( .A0N(N5759), .A1N(n4989), .B0(n6145), .Y(n3745) );
  OAI2BB1X1 U7163 ( .A0N(N5495), .A1N(n5003), .B0(n6296), .Y(n3902) );
  INVX2 U7164 ( .A(reg_length0[3]), .Y(n5956) );
  OAI2BB1X1 U7165 ( .A0N(N5719), .A1N(n4998), .B0(n6193), .Y(n3799) );
  OAI2BB1X1 U7166 ( .A0N(N5715), .A1N(n4998), .B0(n6197), .Y(n3803) );
  OAI2BB1X1 U7167 ( .A0N(N5714), .A1N(n4998), .B0(n6198), .Y(n3804) );
  OAI2BB1X1 U7168 ( .A0N(N5716), .A1N(n4998), .B0(n6196), .Y(n3802) );
  OAI2BB1X1 U7169 ( .A0N(N5717), .A1N(n4998), .B0(n6195), .Y(n3801) );
  OAI2BB1X1 U7170 ( .A0N(N5718), .A1N(n4998), .B0(n6194), .Y(n3800) );
  OAI2BB1X1 U7171 ( .A0N(N5537), .A1N(n5002), .B0(n6244), .Y(n3855) );
  OAI2BB1X1 U7172 ( .A0N(N5800), .A1N(n4991), .B0(n6097), .Y(n3690) );
  OAI2BB1X1 U7173 ( .A0N(N5842), .A1N(n4990), .B0(n6048), .Y(n3634) );
  OAI2BB1X1 U7174 ( .A0N(N5841), .A1N(n4990), .B0(n6049), .Y(n3635) );
  OAI2BB1X1 U7175 ( .A0N(N5534), .A1N(n5002), .B0(n6247), .Y(n3858) );
  OAI2BB1X1 U7176 ( .A0N(N5533), .A1N(n5002), .B0(n6248), .Y(n3859) );
  OAI2BB1X1 U7177 ( .A0N(N5535), .A1N(n5002), .B0(n6246), .Y(n3857) );
  OAI2BB1X1 U7178 ( .A0N(N5536), .A1N(n5002), .B0(n6245), .Y(n3856) );
  OAI2BB1X1 U7179 ( .A0N(N5449), .A1N(n5005), .B0(n5914), .Y(n3947) );
  OAI2BB1X1 U7180 ( .A0N(N5497), .A1N(n5003), .B0(n6294), .Y(n3900) );
  OAI2BB1X1 U7181 ( .A0N(N5496), .A1N(n5003), .B0(n6295), .Y(n3901) );
  OR2X1 U7182 ( .A(n6618), .B(n6661), .Y(n6619) );
  OR2X1 U7183 ( .A(n6613), .B(n6661), .Y(n6614) );
  OAI2BB1X1 U7184 ( .A0N(N5796), .A1N(n4991), .B0(n6101), .Y(n3694) );
  OAI2BB1X1 U7185 ( .A0N(N5448), .A1N(n5005), .B0(n5915), .Y(n3948) );
  OAI2BB1X1 U7186 ( .A0N(N5447), .A1N(n5005), .B0(n5916), .Y(n3949) );
  OAI2BB1X1 U7187 ( .A0N(N5492), .A1N(n5003), .B0(n6299), .Y(n3905) );
  OAI2BB1X1 U7188 ( .A0N(N5493), .A1N(n5003), .B0(n6298), .Y(n3904) );
  OAI2BB1X1 U7189 ( .A0N(N5494), .A1N(n5003), .B0(n6297), .Y(n3903) );
  OAI2BB1X1 U7190 ( .A0N(N5837), .A1N(n4990), .B0(n6053), .Y(n3639) );
  OR2X1 U7191 ( .A(n6569), .B(n6605), .Y(n6570) );
  OAI2BB1X1 U7192 ( .A0N(N5835), .A1N(n4990), .B0(n6055), .Y(n3641) );
  OR2X1 U7193 ( .A(n6674), .B(n6716), .Y(n6675) );
  OR2X1 U7194 ( .A(n6669), .B(n6716), .Y(n6670) );
  OAI2BB1X1 U7195 ( .A0N(N5839), .A1N(n4990), .B0(n6051), .Y(n3637) );
  OAI2BB1X1 U7196 ( .A0N(N5712), .A1N(n4998), .B0(n6200), .Y(n3806) );
  OR2X1 U7197 ( .A(n6736), .B(n6771), .Y(n6737) );
  OR2X1 U7198 ( .A(n6507), .B(n6549), .Y(n6508) );
  OR2X1 U7199 ( .A(n6502), .B(n6549), .Y(n6503) );
  OR2X1 U7200 ( .A(n6557), .B(n6605), .Y(n6558) );
  OR2X1 U7201 ( .A(n6563), .B(n6605), .Y(n6564) );
  OR2X1 U7202 ( .A(n6559), .B(n6605), .Y(n6560) );
  OAI2BB1X1 U7203 ( .A0N(N5838), .A1N(n4990), .B0(n6052), .Y(n3638) );
  OR2X1 U7204 ( .A(n6400), .B(n6441), .Y(n6401) );
  OR2X1 U7205 ( .A(n6395), .B(n6441), .Y(n6396) );
  OR2X1 U7206 ( .A(n6346), .B(n6387), .Y(n6347) );
  OR2X1 U7207 ( .A(n6341), .B(n6387), .Y(n6342) );
  OAI2BB1X1 U7208 ( .A0N(N5531), .A1N(n5002), .B0(n6250), .Y(n3861) );
  OAI2BB1X1 U7209 ( .A0N(N5834), .A1N(n4990), .B0(n6056), .Y(n3642) );
  OAI2BB1X1 U7210 ( .A0N(N5833), .A1N(n4990), .B0(n6057), .Y(n3643) );
  OAI2BB1X1 U7211 ( .A0N(N5799), .A1N(n4991), .B0(n6098), .Y(n3691) );
  OAI2BB1X1 U7212 ( .A0N(N5797), .A1N(n4991), .B0(n6100), .Y(n3693) );
  OAI2BB1X1 U7213 ( .A0N(N5798), .A1N(n4991), .B0(n6099), .Y(n3692) );
  OR2X1 U7214 ( .A(n6513), .B(n6549), .Y(n6514) );
  OAI2BB1X1 U7215 ( .A0N(N5450), .A1N(n5005), .B0(n5913), .Y(n3946) );
  OAI2BB1X1 U7216 ( .A0N(N5710), .A1N(n4998), .B0(n6202), .Y(n3808) );
  OAI2BB1X1 U7217 ( .A0N(N5532), .A1N(n5002), .B0(n6249), .Y(n3860) );
  INVX2 U7218 ( .A(x_in7[0]), .Y(n5468) );
  OR2X1 U7219 ( .A(n6454), .B(n6495), .Y(n6455) );
  OR2X1 U7220 ( .A(n6449), .B(n6495), .Y(n6450) );
  OAI2BB1X1 U7221 ( .A0N(N5752), .A1N(n4989), .B0(n6152), .Y(n3752) );
  OAI2BB1X1 U7222 ( .A0N(N5490), .A1N(n5003), .B0(n6301), .Y(n3907) );
  OAI2BB1X1 U7223 ( .A0N(N5530), .A1N(n5002), .B0(n6251), .Y(n3862) );
  OAI2BB1X1 U7224 ( .A0N(N5529), .A1N(n5002), .B0(n6252), .Y(n3863) );
  OAI221X1 U7225 ( .A0(n6031), .A1(n6039), .B0(n6037), .B1(n6032), .C0(n6783), 
        .Y(n3990) );
  INVX2 U7226 ( .A(reg_length0[4]), .Y(n6031) );
  OAI2BB1X1 U7227 ( .A0N(N5489), .A1N(n5003), .B0(n6302), .Y(n3908) );
  OAI2BB1X1 U7228 ( .A0N(N5488), .A1N(n5003), .B0(n6303), .Y(n3909) );
  OAI2BB1X1 U7229 ( .A0N(N5836), .A1N(n4990), .B0(n6054), .Y(n3640) );
  OR2X1 U7230 ( .A(n6725), .B(n6771), .Y(n6726) );
  OAI2BB1X1 U7231 ( .A0N(N5755), .A1N(n4989), .B0(n6149), .Y(n3749) );
  OAI2BB1X1 U7232 ( .A0N(N5756), .A1N(n4989), .B0(n6148), .Y(n3748) );
  OAI2BB1X1 U7233 ( .A0N(N5757), .A1N(n4989), .B0(n6147), .Y(n3747) );
  OR2X1 U7234 ( .A(n6730), .B(n6771), .Y(n6731) );
  OAI2BB1X1 U7235 ( .A0N(N5713), .A1N(n4998), .B0(n6199), .Y(n3805) );
  OR2X1 U7236 ( .A(n6565), .B(n6605), .Y(n6566) );
  OAI2BB1X1 U7237 ( .A0N(N5491), .A1N(n5003), .B0(n6300), .Y(n3906) );
  OR2X1 U7238 ( .A(n6620), .B(n6661), .Y(n6621) );
  OAI2BB1X1 U7239 ( .A0N(N6365), .A1N(n4999), .B0(n6510), .Y(n3365) );
  OR2X1 U7240 ( .A(n6509), .B(n6549), .Y(n6510) );
  OAI221X1 U7241 ( .A0(n6039), .A1(n6038), .B0(n6037), .B1(n6040), .C0(n6782), 
        .Y(n4028) );
  INVX2 U7242 ( .A(reg_length0[5]), .Y(n6038) );
  OAI2BB1X1 U7243 ( .A0N(N5753), .A1N(n4989), .B0(n6151), .Y(n3751) );
  OR2X1 U7244 ( .A(n6402), .B(n6441), .Y(n6403) );
  OR2X1 U7245 ( .A(n6348), .B(n6387), .Y(n6349) );
  OAI2BB1X1 U7246 ( .A0N(N5793), .A1N(n4991), .B0(n6104), .Y(n3697) );
  OAI2BB1X1 U7247 ( .A0N(N5792), .A1N(n4991), .B0(n6105), .Y(n3698) );
  OR2X1 U7248 ( .A(n6676), .B(n6716), .Y(n6677) );
  OAI2BB1X1 U7249 ( .A0N(N5751), .A1N(n4989), .B0(n6153), .Y(n3753) );
  OR2X1 U7250 ( .A(n6680), .B(n6716), .Y(n6681) );
  OR2X1 U7251 ( .A(n6352), .B(n6387), .Y(n6353) );
  OAI2BB1XL U7252 ( .A0N(reg_length00[5]), .A1N(n6787), .B0(n6782), .Y(n3171)
         );
  OAI2BB1XL U7253 ( .A0N(reg_length00[4]), .A1N(n6787), .B0(n6783), .Y(n3172)
         );
  OR2X1 U7254 ( .A(n6732), .B(n6771), .Y(n6733) );
  OR2X1 U7255 ( .A(n6406), .B(n6441), .Y(n6407) );
  OAI2BB1X1 U7256 ( .A0N(N5709), .A1N(n4998), .B0(n6203), .Y(n3809) );
  OAI2BB1X1 U7257 ( .A0N(N5754), .A1N(n4989), .B0(n6150), .Y(n3750) );
  OR2X1 U7258 ( .A(n6460), .B(n6495), .Y(n6461) );
  OR2X1 U7259 ( .A(n6624), .B(n6661), .Y(n6625) );
  OR2X1 U7260 ( .A(n6456), .B(n6495), .Y(n6457) );
  OAI2BB1X1 U7261 ( .A0N(N5794), .A1N(n4991), .B0(n6103), .Y(n3696) );
  NAND2X1 U7262 ( .A(n5973), .B(n6779), .Y(n3991) );
  MXI2X1 U7263 ( .A(n5958), .B(n5957), .S0(reg_length0[0]), .Y(n5973) );
  INVX2 U7264 ( .A(n6039), .Y(n5957) );
  OAI2BB1X1 U7265 ( .A0N(N5707), .A1N(n4998), .B0(n6205), .Y(n3811) );
  OAI2BB1X1 U7266 ( .A0N(N5708), .A1N(n4998), .B0(n6204), .Y(n3810) );
  OAI2BB1X1 U7267 ( .A0N(N5485), .A1N(n5003), .B0(n6306), .Y(n3912) );
  OAI2BB1X1 U7268 ( .A0N(N5486), .A1N(n5003), .B0(n6305), .Y(n3911) );
  OAI221X1 U7269 ( .A0(n6025), .A1(n6039), .B0(n5344), .B1(n6037), .C0(n6785), 
        .Y(n3988) );
  INVX2 U7270 ( .A(reg_length0[2]), .Y(n6025) );
  OAI2BB1X1 U7271 ( .A0N(N5446), .A1N(n5005), .B0(n5917), .Y(n3950) );
  OR2X1 U7272 ( .A(n4958), .B(n6605), .Y(n6571) );
  OR2X1 U7273 ( .A(n4959), .B(n6771), .Y(n6738) );
  OAI2BB1X1 U7274 ( .A0N(N5832), .A1N(n4990), .B0(n6058), .Y(n3644) );
  OR2X1 U7275 ( .A(n4960), .B(n6549), .Y(n6515) );
  OAI2BB1X1 U7276 ( .A0N(N5528), .A1N(n5002), .B0(n6253), .Y(n3864) );
  OR2X1 U7277 ( .A(n6682), .B(n6716), .Y(n6683) );
  OAI2BB1X1 U7278 ( .A0N(N5487), .A1N(n5003), .B0(n6304), .Y(n3910) );
  OAI2BB1X1 U7279 ( .A0N(N5706), .A1N(n4998), .B0(n6206), .Y(n3812) );
  OAI2BB1X1 U7280 ( .A0N(N5484), .A1N(n5003), .B0(n6307), .Y(n3913) );
  OAI2BB1X1 U7281 ( .A0N(N5444), .A1N(n5005), .B0(n5919), .Y(n3952) );
  OAI2BB1X1 U7282 ( .A0N(N5445), .A1N(n5005), .B0(n5918), .Y(n3951) );
  OAI2BB1X1 U7283 ( .A0N(N5791), .A1N(n4991), .B0(n6106), .Y(n3699) );
  OAI2BB1X1 U7284 ( .A0N(N5526), .A1N(n5002), .B0(n6255), .Y(n3866) );
  OAI2BB1X1 U7285 ( .A0N(N5527), .A1N(n5002), .B0(n6254), .Y(n3865) );
  OAI2BB1X1 U7286 ( .A0N(N5750), .A1N(n4989), .B0(n6154), .Y(n3754) );
  OR2X1 U7287 ( .A(n6354), .B(n6387), .Y(n6355) );
  OAI2BB1X1 U7288 ( .A0N(N5831), .A1N(n4990), .B0(n6059), .Y(n3645) );
  OR2X1 U7289 ( .A(n6408), .B(n6441), .Y(n6409) );
  OR2X1 U7290 ( .A(n6686), .B(n6716), .Y(n6687) );
  OAI2BB1X1 U7291 ( .A0N(N5830), .A1N(n4990), .B0(n6060), .Y(n3646) );
  OR2X1 U7292 ( .A(n6462), .B(n6495), .Y(n6463) );
  OR2X1 U7293 ( .A(n6626), .B(n6661), .Y(n6627) );
  OAI2BB1X1 U7294 ( .A0N(N5748), .A1N(n4989), .B0(n6156), .Y(n3756) );
  OAI2BB1X1 U7295 ( .A0N(N5749), .A1N(n4989), .B0(n6155), .Y(n3755) );
  OAI2BB1X1 U7296 ( .A0N(N5789), .A1N(n4991), .B0(n6108), .Y(n3701) );
  OAI2BB1X1 U7297 ( .A0N(N5790), .A1N(n4991), .B0(n6107), .Y(n3700) );
  OR2X1 U7298 ( .A(n4955), .B(n6441), .Y(n6412) );
  OR2X1 U7299 ( .A(n6574), .B(n6605), .Y(n6575) );
  OAI2BB1X1 U7300 ( .A0N(N5443), .A1N(n5005), .B0(n5920), .Y(n3953) );
  OR2X1 U7301 ( .A(n6741), .B(n6771), .Y(n6742) );
  OR2X1 U7302 ( .A(n6630), .B(n6661), .Y(n6631) );
  OAI2BB1X1 U7303 ( .A0N(N5829), .A1N(n4990), .B0(n6061), .Y(n3647) );
  OR2X1 U7304 ( .A(n4961), .B(n6771), .Y(n6743) );
  OAI2BB1X1 U7305 ( .A0N(N5828), .A1N(n4990), .B0(n6062), .Y(n3648) );
  OR2X1 U7306 ( .A(n6518), .B(n6549), .Y(n6519) );
  OAI2BB1X1 U7307 ( .A0N(N5525), .A1N(n5002), .B0(n6256), .Y(n3867) );
  OAI2BB1X1 U7308 ( .A0N(N5524), .A1N(n5002), .B0(n6257), .Y(n3868) );
  OR2X1 U7309 ( .A(n4956), .B(n6495), .Y(n6466) );
  OAI2BB1X1 U7310 ( .A0N(N5705), .A1N(n4998), .B0(n6207), .Y(n3813) );
  OAI2BB1X1 U7311 ( .A0N(N5788), .A1N(n4991), .B0(n6109), .Y(n3702) );
  OAI2BB1X1 U7312 ( .A0N(N5787), .A1N(n4991), .B0(n6110), .Y(n3703) );
  OAI2BB1X1 U7313 ( .A0N(N5747), .A1N(n4989), .B0(n6157), .Y(n3757) );
  OR2X1 U7314 ( .A(n4957), .B(n6387), .Y(n6358) );
  OR2X1 U7315 ( .A(n4962), .B(n6387), .Y(n6359) );
  OAI2BB1X1 U7316 ( .A0N(N5746), .A1N(n4989), .B0(n6158), .Y(n3758) );
  OR2X1 U7317 ( .A(n6576), .B(n6605), .Y(n6577) );
  OAI2BB1X1 U7318 ( .A0N(N5442), .A1N(n5005), .B0(n5921), .Y(n3954) );
  OR2X1 U7319 ( .A(n4963), .B(n6495), .Y(n6467) );
  OAI2BB1X1 U7320 ( .A0N(N5483), .A1N(n5003), .B0(n6308), .Y(n3914) );
  OR2X1 U7321 ( .A(n6520), .B(n6549), .Y(n6521) );
  OR2X1 U7322 ( .A(n4964), .B(n6716), .Y(n6688) );
  OR2X1 U7323 ( .A(n4965), .B(n6441), .Y(n6413) );
  OAI2BB1X1 U7324 ( .A0N(N5826), .A1N(n4990), .B0(n6064), .Y(n3650) );
  OAI2BB1X1 U7325 ( .A0N(N5480), .A1N(n5003), .B0(n6312), .Y(n3917) );
  OR2X1 U7326 ( .A(n6336), .B(n6311), .Y(n6312) );
  INVX2 U7327 ( .A(y_out_sum1[19]), .Y(n6311) );
  OAI2BB1X1 U7328 ( .A0N(N5522), .A1N(n5002), .B0(n6259), .Y(n3870) );
  OAI2BB1X1 U7329 ( .A0N(N5523), .A1N(n5002), .B0(n6258), .Y(n3869) );
  OAI2BB1X1 U7330 ( .A0N(N6275), .A1N(n4996), .B0(n6633), .Y(n3483) );
  OR2X1 U7331 ( .A(n6632), .B(n6661), .Y(n6633) );
  OAI2BB1X1 U7332 ( .A0N(N5482), .A1N(n5003), .B0(n6309), .Y(n3915) );
  OAI2BB1X1 U7333 ( .A0N(N5827), .A1N(n4990), .B0(n6063), .Y(n3649) );
  OAI2BB1X1 U7334 ( .A0N(N5786), .A1N(n4991), .B0(n6111), .Y(n3704) );
  OAI2BB1X1 U7335 ( .A0N(N5744), .A1N(n4989), .B0(n6160), .Y(n3760) );
  OAI2BB1X1 U7336 ( .A0N(N5703), .A1N(n4998), .B0(n6209), .Y(n3815) );
  OAI2BB1X1 U7337 ( .A0N(N5745), .A1N(n4989), .B0(n6159), .Y(n3759) );
  OAI2BB1X1 U7338 ( .A0N(N5441), .A1N(n5005), .B0(n5922), .Y(n3955) );
  OAI2BB1X1 U7339 ( .A0N(N5704), .A1N(n4998), .B0(n6208), .Y(n3814) );
  OAI2BB1X1 U7340 ( .A0N(N5825), .A1N(n4990), .B0(n6066), .Y(n3651) );
  OR2X1 U7341 ( .A(n6090), .B(n6065), .Y(n6066) );
  INVX2 U7342 ( .A(y_out_sum6[19]), .Y(n6065) );
  OAI2BB1X1 U7343 ( .A0N(N5743), .A1N(n4989), .B0(n6162), .Y(n3761) );
  OR2X1 U7344 ( .A(n6186), .B(n6161), .Y(n6162) );
  INVX2 U7345 ( .A(y_out_sum4[19]), .Y(n6161) );
  OAI2BB1X1 U7346 ( .A0N(N5481), .A1N(n5003), .B0(n6310), .Y(n3916) );
  OAI2BB1X1 U7347 ( .A0N(N5785), .A1N(n4991), .B0(n6112), .Y(n3705) );
  OAI2BB1X1 U7348 ( .A0N(N5440), .A1N(n5005), .B0(n5923), .Y(n3956) );
  OAI2BB1X1 U7349 ( .A0N(N5824), .A1N(n4990), .B0(n6068), .Y(n3652) );
  OR2X1 U7350 ( .A(n6090), .B(n6067), .Y(n6068) );
  INVX2 U7351 ( .A(y_out_sum6[18]), .Y(n6067) );
  OAI2BB1X1 U7352 ( .A0N(N5699), .A1N(n4998), .B0(n6216), .Y(n3819) );
  OR2X1 U7353 ( .A(n6235), .B(n6215), .Y(n6216) );
  INVX2 U7354 ( .A(y_out_sum3[16]), .Y(n6215) );
  NAND3X1 U7355 ( .A(in_valid), .B(n117), .C(n1312), .Y(n2732) );
  AND4X2 U7356 ( .A(n2625), .B(n2626), .C(n2627), .D(n2628), .Y(n2624) );
  AOI222XL U7357 ( .A0(N5059), .A1(n2568), .B0(N5067), .B1(n2559), .C0(N5075), 
        .C1(n2567), .Y(n2628) );
  AOI221XL U7358 ( .A0(n2560), .A1(count28[1]), .B0(n7233), .B1(w_mat_idx), 
        .C0(n2603), .Y(n2625) );
  AOI222XL U7359 ( .A0(n7172), .A1(count48[1]), .B0(n7171), .B1(count58[1]), 
        .C0(n7173), .C1(count38[1]), .Y(n2626) );
  AOI222XL U7360 ( .A0(n2570), .A1(count78[1]), .B0(n5372), .B1(n2566), .C0(
        n2569), .C1(count68[1]), .Y(n2627) );
  AND4X2 U7361 ( .A(n2643), .B(n2644), .C(n2645), .D(n2646), .Y(n2642) );
  AOI222XL U7362 ( .A0(n7311), .A1(n2567), .B0(n5573), .B1(n2558), .C0(n7311), 
        .C1(n2559), .Y(n2646) );
  AOI221XL U7363 ( .A0(n7172), .A1(count48[0]), .B0(n2560), .B1(count28[0]), 
        .C0(n2603), .Y(n2643) );
  AOI222XL U7364 ( .A0(n2569), .A1(count68[0]), .B0(n5379), .B1(n2568), .C0(
        n5366), .C1(n2566), .Y(n2645) );
  AOI222XL U7365 ( .A0(n7173), .A1(count38[0]), .B0(n2570), .B1(count78[0]), 
        .C0(n7171), .C1(count58[0]), .Y(n2644) );
  OAI2BB1X1 U7366 ( .A0N(N5742), .A1N(n4989), .B0(n6164), .Y(n3762) );
  OR2X1 U7367 ( .A(n6186), .B(n6163), .Y(n6164) );
  INVX2 U7368 ( .A(y_out_sum4[18]), .Y(n6163) );
  OAI2BB1X1 U7369 ( .A0N(N5439), .A1N(n5005), .B0(n5925), .Y(n3957) );
  OR2X1 U7370 ( .A(n5949), .B(n5924), .Y(n5925) );
  INVX2 U7371 ( .A(y_out_sum0[19]), .Y(n5924) );
  OAI2BB1X1 U7372 ( .A0N(N5479), .A1N(n5003), .B0(n6314), .Y(n3918) );
  OR2X1 U7373 ( .A(n6336), .B(n6313), .Y(n6314) );
  INVX2 U7374 ( .A(y_out_sum1[18]), .Y(n6313) );
  OAI2BB1X1 U7375 ( .A0N(N5521), .A1N(n5002), .B0(n6261), .Y(n3871) );
  OR2X1 U7376 ( .A(n6286), .B(n6260), .Y(n6261) );
  INVX2 U7377 ( .A(y_out_sum2[19]), .Y(n6260) );
  OAI2BB1X1 U7378 ( .A0N(N5784), .A1N(n4991), .B0(n6114), .Y(n3706) );
  OR2X1 U7379 ( .A(n6138), .B(n6113), .Y(n6114) );
  INVX2 U7380 ( .A(y_out_sum5[19]), .Y(n6113) );
  AOI222XL U7381 ( .A0(n7173), .A1(count38[2]), .B0(n2570), .B1(count78[2]), 
        .C0(n7171), .C1(count58[2]), .Y(n2608) );
  OR2X1 U7382 ( .A(n2605), .B(n2606), .Y(N5147) );
  NAND4X1 U7383 ( .A(n2615), .B(n2616), .C(n2617), .D(n2618), .Y(n2605) );
  NAND4X1 U7384 ( .A(n2607), .B(n2608), .C(n2609), .D(n2610), .Y(n2606) );
  AOI221XL U7385 ( .A0(temp_w_mat_idx[0]), .A1(n2591), .B0(n7030), .B1(n2619), 
        .C0(n2620), .Y(n2618) );
  OAI2BB1X1 U7386 ( .A0N(N5702), .A1N(n4998), .B0(n6211), .Y(n3816) );
  OR2X1 U7387 ( .A(n6235), .B(n6210), .Y(n6211) );
  INVX2 U7388 ( .A(y_out_sum3[19]), .Y(n6210) );
  OAI2BB1X1 U7389 ( .A0N(N5698), .A1N(n4998), .B0(n6218), .Y(n3820) );
  OR2X1 U7390 ( .A(n6235), .B(n6217), .Y(n6218) );
  INVX2 U7391 ( .A(y_out_sum3[15]), .Y(n6217) );
  OAI2BB1X1 U7392 ( .A0N(N5520), .A1N(n5002), .B0(n6263), .Y(n3872) );
  OR2X1 U7393 ( .A(n6286), .B(n6262), .Y(n6263) );
  INVX2 U7394 ( .A(y_out_sum2[18]), .Y(n6262) );
  OAI2BB1X1 U7395 ( .A0N(N5701), .A1N(n4998), .B0(n6213), .Y(n3817) );
  OR2X1 U7396 ( .A(n6235), .B(n6212), .Y(n6213) );
  INVX2 U7397 ( .A(y_out_sum3[18]), .Y(n6212) );
  OAI2BB1X1 U7398 ( .A0N(N5438), .A1N(n5005), .B0(n5927), .Y(n3958) );
  OR2X1 U7399 ( .A(n5949), .B(n5926), .Y(n5927) );
  INVX2 U7400 ( .A(y_out_sum0[18]), .Y(n5926) );
  AOI222XL U7401 ( .A0(n2569), .A1(count68[2]), .B0(n5571), .B1(n2568), .C0(
        n5371), .C1(n2566), .Y(n2609) );
  OAI2BB1X1 U7402 ( .A0N(N6229), .A1N(n4995), .B0(n6693), .Y(n3543) );
  OAI2BB1X1 U7403 ( .A0N(N5823), .A1N(n4990), .B0(n6069), .Y(n3653) );
  OAI2BB1X1 U7404 ( .A0N(N6311), .A1N(n4997), .B0(n6582), .Y(n3433) );
  OAI2BB1X1 U7405 ( .A0N(N5783), .A1N(n4991), .B0(n6116), .Y(n3707) );
  OR2X1 U7406 ( .A(n6138), .B(n6115), .Y(n6116) );
  INVX2 U7407 ( .A(y_out_sum5[18]), .Y(n6115) );
  OAI2BB1X1 U7408 ( .A0N(N6188), .A1N(n4994), .B0(n6748), .Y(n3598) );
  NAND4X1 U7409 ( .A(n2540), .B(n2541), .C(n2542), .D(n2543), .Y(N5151) );
  AND4X2 U7410 ( .A(n2544), .B(n2545), .C(n2546), .D(n2547), .Y(n2543) );
  AOI222XL U7411 ( .A0(n5367), .A1(n2566), .B0(N5080), .B1(n2567), .C0(N5064), 
        .C1(n2568), .Y(n2541) );
  AOI22X1 U7412 ( .A0(n2569), .A1(count68[6]), .B0(n2570), .B1(count78[6]), 
        .Y(n2540) );
  NAND4X1 U7413 ( .A(n2571), .B(n2572), .C(n2573), .D(n2574), .Y(N5150) );
  AOI222XL U7414 ( .A0(n5567), .A1(n2568), .B0(N5071), .B1(n2559), .C0(N5079), 
        .C1(n2567), .Y(n2572) );
  AND4X2 U7415 ( .A(n2575), .B(n2576), .C(n2577), .D(n2578), .Y(n2574) );
  AOI222XL U7416 ( .A0(n2570), .A1(count78[5]), .B0(n5368), .B1(n2566), .C0(
        n2569), .C1(count68[5]), .Y(n2571) );
  NAND4X1 U7417 ( .A(n2582), .B(n2583), .C(n2584), .D(n2585), .Y(N5149) );
  AOI222XL U7418 ( .A0(n5568), .A1(n2568), .B0(N5070), .B1(n2559), .C0(N5078), 
        .C1(n2567), .Y(n2583) );
  AND4X2 U7419 ( .A(n2586), .B(n2587), .C(n2588), .D(n2589), .Y(n2585) );
  AOI222XL U7420 ( .A0(n2570), .A1(count78[4]), .B0(n5369), .B1(n2566), .C0(
        n2569), .C1(count68[4]), .Y(n2582) );
  NAND4X1 U7421 ( .A(n2593), .B(n2594), .C(n2595), .D(n2596), .Y(N5148) );
  AOI222XL U7422 ( .A0(N5061), .A1(n2568), .B0(N5069), .B1(n2559), .C0(N5077), 
        .C1(n2567), .Y(n2594) );
  AND4X2 U7423 ( .A(n2597), .B(n2598), .C(n2599), .D(n2600), .Y(n2596) );
  AOI222XL U7424 ( .A0(n2570), .A1(count78[3]), .B0(n5370), .B1(n2566), .C0(
        n2569), .C1(count68[3]), .Y(n2593) );
  AOI221XL U7425 ( .A0(n2560), .A1(count28[3]), .B0(n7231), .B1(w_mat_idx), 
        .C0(n2604), .Y(n2595) );
  OAI222X1 U7426 ( .A0(n7462), .A1(n2563), .B0(n7476), .B1(n2564), .C0(n7469), 
        .C1(n2565), .Y(n2604) );
  AOI221XL U7427 ( .A0(n2560), .A1(count28[5]), .B0(n7231), .B1(
        temp_w_mat_idx[1]), .C0(n2581), .Y(n2573) );
  OAI222X1 U7428 ( .A0(n7464), .A1(n2563), .B0(n7478), .B1(n2564), .C0(n7471), 
        .C1(n2565), .Y(n2581) );
  AOI221XL U7429 ( .A0(n2560), .A1(count28[4]), .B0(n7231), .B1(
        temp_w_mat_idx[0]), .C0(n2592), .Y(n2584) );
  OAI222X1 U7430 ( .A0(n7463), .A1(n2563), .B0(n7477), .B1(n2564), .C0(n7470), 
        .C1(n2565), .Y(n2592) );
  AOI221XL U7431 ( .A0(n2560), .A1(count28[6]), .B0(n7231), .B1(
        temp_w_mat_idx[2]), .C0(n2562), .Y(n2542) );
  OAI222X1 U7432 ( .A0(n7465), .A1(n2563), .B0(n7479), .B1(n2564), .C0(n7472), 
        .C1(n2565), .Y(n2562) );
  OAI2BB1X1 U7433 ( .A0N(N6433), .A1N(n4992), .B0(n6420), .Y(n3269) );
  OR2X1 U7434 ( .A(n6441), .B(n6419), .Y(n6420) );
  INVX2 U7435 ( .A(y_out_sum13[16]), .Y(n6419) );
  OAI2BB1X1 U7436 ( .A0N(N5700), .A1N(n4998), .B0(n6214), .Y(n3818) );
  OAI2BB1X1 U7437 ( .A0N(N5741), .A1N(n4989), .B0(n6165), .Y(n3763) );
  OAI2BB1X1 U7438 ( .A0N(N5478), .A1N(n5003), .B0(n6315), .Y(n3919) );
  OAI2BB1X1 U7439 ( .A0N(N5519), .A1N(n5002), .B0(n6264), .Y(n3873) );
  OAI2BB1X1 U7440 ( .A0N(N5782), .A1N(n4991), .B0(n6117), .Y(n3708) );
  OAI2BB1X1 U7441 ( .A0N(N6352), .A1N(n4999), .B0(n6526), .Y(n3378) );
  OAI2BB1X1 U7442 ( .A0N(N6270), .A1N(n4996), .B0(n6638), .Y(n3488) );
  OAI2BB1X1 U7443 ( .A0N(N5437), .A1N(n5005), .B0(n5928), .Y(n3959) );
  OAI2BB1X1 U7444 ( .A0N(N5477), .A1N(n5003), .B0(n6317), .Y(n3920) );
  OR2X1 U7445 ( .A(n6336), .B(n6316), .Y(n6317) );
  INVX2 U7446 ( .A(y_out_sum1[16]), .Y(n6316) );
  OAI2BB1X1 U7447 ( .A0N(N6392), .A1N(n5000), .B0(n6474), .Y(n3324) );
  OR2X1 U7448 ( .A(n6495), .B(n6473), .Y(n6474) );
  INVX2 U7449 ( .A(y_out_sum12[16]), .Y(n6473) );
  OAI2BB1X1 U7450 ( .A0N(N6187), .A1N(n4994), .B0(n6750), .Y(n3599) );
  OR2X1 U7451 ( .A(n6771), .B(n6749), .Y(n6750) );
  INVX2 U7452 ( .A(y_out_sum7[16]), .Y(n6749) );
  OAI2BB1X1 U7453 ( .A0N(N6393), .A1N(n5000), .B0(n6472), .Y(n3323) );
  OAI2BB1X1 U7454 ( .A0N(N6475), .A1N(n4993), .B0(n6364), .Y(n3213) );
  OAI2BB1X1 U7455 ( .A0N(N5518), .A1N(n5002), .B0(n6266), .Y(n3874) );
  OR2X1 U7456 ( .A(n6286), .B(n6265), .Y(n6266) );
  INVX2 U7457 ( .A(y_out_sum2[16]), .Y(n6265) );
  OAI2BB1X1 U7458 ( .A0N(N6269), .A1N(n4996), .B0(n6640), .Y(n3489) );
  OR2X1 U7459 ( .A(n6661), .B(n6639), .Y(n6640) );
  INVX2 U7460 ( .A(y_out_sum9[16]), .Y(n6639) );
  OAI2BB1X1 U7461 ( .A0N(N6351), .A1N(n4999), .B0(n6528), .Y(n3379) );
  OR2X1 U7462 ( .A(n6549), .B(n6527), .Y(n6528) );
  INVX2 U7463 ( .A(y_out_sum11[16]), .Y(n6527) );
  OAI2BB1X1 U7464 ( .A0N(N6434), .A1N(n4992), .B0(n6418), .Y(n3268) );
  OAI2BB1X1 U7465 ( .A0N(N6310), .A1N(n4997), .B0(n6584), .Y(n3434) );
  OR2X1 U7466 ( .A(n6605), .B(n6583), .Y(n6584) );
  INVX2 U7467 ( .A(y_out_sum10[16]), .Y(n6583) );
  OAI2BB1X1 U7468 ( .A0N(N6228), .A1N(n4995), .B0(n6695), .Y(n3544) );
  OR2X1 U7469 ( .A(n6716), .B(n6694), .Y(n6695) );
  INVX2 U7470 ( .A(y_out_sum8[16]), .Y(n6694) );
  OAI2BB1X1 U7471 ( .A0N(N5781), .A1N(n4991), .B0(n6119), .Y(n3709) );
  OR2X1 U7472 ( .A(n6138), .B(n6118), .Y(n6119) );
  INVX2 U7473 ( .A(y_out_sum5[16]), .Y(n6118) );
  OAI2BB1X1 U7474 ( .A0N(N5436), .A1N(n5005), .B0(n5930), .Y(n3960) );
  OR2X1 U7475 ( .A(n5949), .B(n5929), .Y(n5930) );
  INVX2 U7476 ( .A(y_out_sum0[16]), .Y(n5929) );
  OAI2BB1X1 U7477 ( .A0N(N5476), .A1N(n5003), .B0(n6319), .Y(n3921) );
  OR2X1 U7478 ( .A(n6336), .B(n6318), .Y(n6319) );
  INVX2 U7479 ( .A(y_out_sum1[15]), .Y(n6318) );
  OAI2BB1X1 U7480 ( .A0N(N6474), .A1N(n4993), .B0(n6366), .Y(n3214) );
  OR2X1 U7481 ( .A(n6387), .B(n6365), .Y(n6366) );
  INVX2 U7482 ( .A(y_out_sum14[16]), .Y(n6365) );
  OAI2BB1X1 U7483 ( .A0N(N5822), .A1N(n4990), .B0(n6071), .Y(n3654) );
  OR2X1 U7484 ( .A(n6090), .B(n6070), .Y(n6071) );
  INVX2 U7485 ( .A(y_out_sum6[16]), .Y(n6070) );
  OAI2BB1X1 U7486 ( .A0N(N5740), .A1N(n4989), .B0(n6167), .Y(n3764) );
  OR2X1 U7487 ( .A(n6186), .B(n6166), .Y(n6167) );
  INVX2 U7488 ( .A(y_out_sum4[16]), .Y(n6166) );
  OAI2BB1X1 U7489 ( .A0N(N5517), .A1N(n5002), .B0(n6268), .Y(n3875) );
  OR2X1 U7490 ( .A(n6286), .B(n6267), .Y(n6268) );
  INVX2 U7491 ( .A(y_out_sum2[15]), .Y(n6267) );
  OAI2BB1X1 U7492 ( .A0N(N5697), .A1N(n4998), .B0(n6219), .Y(n3821) );
  OAI2BB1X1 U7493 ( .A0N(N5821), .A1N(n4990), .B0(n6073), .Y(n3655) );
  OR2X1 U7494 ( .A(n6090), .B(n6072), .Y(n6073) );
  INVX2 U7495 ( .A(y_out_sum6[15]), .Y(n6072) );
  NAND3X1 U7496 ( .A(in_valid), .B(n5465), .C(n1312), .Y(n2671) );
  OAI2BB1X1 U7497 ( .A0N(N5780), .A1N(n4991), .B0(n6121), .Y(n3710) );
  OR2X1 U7498 ( .A(n6138), .B(n6120), .Y(n6121) );
  INVX2 U7499 ( .A(y_out_sum5[15]), .Y(n6120) );
  OAI2BB1X1 U7500 ( .A0N(N5435), .A1N(n5005), .B0(n5932), .Y(n3961) );
  OR2X1 U7501 ( .A(n5949), .B(n5931), .Y(n5932) );
  INVX2 U7502 ( .A(y_out_sum0[15]), .Y(n5931) );
  OAI2BB1X1 U7503 ( .A0N(N5475), .A1N(n5003), .B0(n6320), .Y(n3922) );
  OAI2BB1X1 U7504 ( .A0N(N5738), .A1N(n4989), .B0(n6170), .Y(n3766) );
  OAI2BB1X1 U7505 ( .A0N(N5434), .A1N(n5005), .B0(n5933), .Y(n3962) );
  OAI2BB1X1 U7506 ( .A0N(N5739), .A1N(n4989), .B0(n6169), .Y(n3765) );
  OR2X1 U7507 ( .A(n6186), .B(n6168), .Y(n6169) );
  INVX2 U7508 ( .A(y_out_sum4[15]), .Y(n6168) );
  AOI222XL U7509 ( .A0(n7208), .A1(w_mat_idx), .B0(n7172), .B1(count48[2]), 
        .C0(n2560), .C1(count28[2]), .Y(n2607) );
  OAI2BB1X1 U7510 ( .A0N(N5516), .A1N(n5002), .B0(n6269), .Y(n3876) );
  OAI2BB1X1 U7511 ( .A0N(N5779), .A1N(n4991), .B0(n6122), .Y(n3711) );
  OAI2BB1X1 U7512 ( .A0N(N5820), .A1N(n4990), .B0(n6074), .Y(n3656) );
  OAI2BB1X1 U7513 ( .A0N(N5819), .A1N(n4990), .B0(n6075), .Y(n3657) );
  OAI2BB1X1 U7514 ( .A0N(N6266), .A1N(n4996), .B0(n6643), .Y(n3492) );
  AOI222XL U7515 ( .A0(N5139), .A1(n2553), .B0(n7176), .B1(count08[1]), .C0(
        n7174), .C1(count18[1]), .Y(n2633) );
  AOI222XL U7516 ( .A0(N5142), .A1(n2553), .B0(n7176), .B1(count08[4]), .C0(
        n7174), .C1(count18[4]), .Y(n2588) );
  AOI222XL U7517 ( .A0(N5141), .A1(n2553), .B0(n7176), .B1(count08[3]), .C0(
        n7174), .C1(count18[3]), .Y(n2599) );
  OAI2BB1X1 U7518 ( .A0N(N6225), .A1N(n4995), .B0(n6698), .Y(n3547) );
  AOI222XL U7519 ( .A0(N5127), .A1(n2554), .B0(n7174), .B1(count18[5]), .C0(
        N5143), .C1(n2553), .Y(n2577) );
  OAI2BB1X1 U7520 ( .A0N(N6184), .A1N(n4994), .B0(n6753), .Y(n3602) );
  OAI2BB1X1 U7521 ( .A0N(N5818), .A1N(n4990), .B0(n6076), .Y(n3658) );
  AOI222XL U7522 ( .A0(n7174), .A1(count18[6]), .B0(temp_w_mat_idx[3]), .B1(
        n7229), .C0(n7176), .C1(count08[6]), .Y(n2547) );
  INVX2 U7523 ( .A(n2551), .Y(n7229) );
  OAI2BB1X1 U7524 ( .A0N(N6430), .A1N(n4992), .B0(n6423), .Y(n3272) );
  OAI2BB1X1 U7525 ( .A0N(N6348), .A1N(n4999), .B0(n6531), .Y(n3382) );
  OAI2BB1X1 U7526 ( .A0N(N5474), .A1N(n5003), .B0(n6321), .Y(n3923) );
  OAI2BB1X1 U7527 ( .A0N(N6224), .A1N(n4995), .B0(n6699), .Y(n3548) );
  OAI2BB1X1 U7528 ( .A0N(N6470), .A1N(n4993), .B0(n6370), .Y(n3218) );
  OAI2BB1X1 U7529 ( .A0N(N5736), .A1N(n4989), .B0(n6172), .Y(n3768) );
  AOI222XL U7530 ( .A0(n7174), .A1(count18[2]), .B0(temp_w_mat_idx[1]), .B1(
        n2590), .C0(n7176), .C1(count08[2]), .Y(n2617) );
  OAI2BB1X1 U7531 ( .A0N(N6183), .A1N(n4994), .B0(n6754), .Y(n3603) );
  OAI2BB1X1 U7532 ( .A0N(N6306), .A1N(n4997), .B0(n6588), .Y(n3438) );
  OAI2BB1X1 U7533 ( .A0N(N5737), .A1N(n4989), .B0(n6171), .Y(n3767) );
  OAI2BB1X1 U7534 ( .A0N(N5515), .A1N(n5002), .B0(n6270), .Y(n3877) );
  OAI2BB1X1 U7535 ( .A0N(N6307), .A1N(n4997), .B0(n6587), .Y(n3437) );
  OAI2BB1X1 U7536 ( .A0N(N5433), .A1N(n5005), .B0(n5934), .Y(n3963) );
  OAI2BB1X1 U7537 ( .A0N(N5778), .A1N(n4991), .B0(n6123), .Y(n3712) );
  OAI2BB1X1 U7538 ( .A0N(N6388), .A1N(n5000), .B0(n6478), .Y(n3328) );
  OAI2BB1X1 U7539 ( .A0N(N5696), .A1N(n4998), .B0(n6220), .Y(n3822) );
  OAI2BB1X1 U7540 ( .A0N(N6471), .A1N(n4993), .B0(n6369), .Y(n3217) );
  OAI2BB1X1 U7541 ( .A0N(N5695), .A1N(n4998), .B0(n6221), .Y(n3823) );
  OAI2BB1X1 U7542 ( .A0N(N6389), .A1N(n5000), .B0(n6477), .Y(n3327) );
  AOI222XL U7543 ( .A0(n7176), .A1(count08[5]), .B0(temp_w_mat_idx[2]), .B1(
        n2579), .C0(temp_w_mat_idx[3]), .C1(n2580), .Y(n2578) );
  NOR3X1 U7544 ( .A(reg_invalid2[7]), .B(reg_invalid2[8]), .C(reg_invalid2[6]), 
        .Y(n2715) );
  NAND3X1 U7545 ( .A(reg_invalid2[4]), .B(n2715), .C(n5373), .Y(n2814) );
  NAND4BX1 U7546 ( .AN(n1907), .B(n1585), .C(n2702), .D(n2703), .Y(n2619) );
  AOI22X1 U7547 ( .A0(n2716), .A1(n7044), .B0(n7328), .B1(n2717), .Y(n2702) );
  AOI211X1 U7548 ( .A0(n7046), .A1(reg_invalid2[0]), .B0(n2674), .C0(n2637), 
        .Y(n2703) );
  OAI2BB1X1 U7549 ( .A0N(N5514), .A1N(n5002), .B0(n6271), .Y(n3878) );
  OAI2BB1X1 U7550 ( .A0N(N5777), .A1N(n4991), .B0(n6124), .Y(n3713) );
  OAI2BB1X1 U7551 ( .A0N(N6265), .A1N(n4996), .B0(n6644), .Y(n3493) );
  OAI2BB1X1 U7552 ( .A0N(N5432), .A1N(n5005), .B0(n5935), .Y(n3964) );
  OAI2BB1X1 U7553 ( .A0N(N5735), .A1N(n4989), .B0(n6173), .Y(n3769) );
  NAND2X1 U7554 ( .A(in_valid), .B(n5457), .Y(n1313) );
  NAND2X1 U7555 ( .A(N5006), .B(n7177), .Y(n2670) );
  OAI2BB1X1 U7556 ( .A0N(N5473), .A1N(n5003), .B0(n6322), .Y(n3924) );
  OAI2BB1X1 U7557 ( .A0N(N6347), .A1N(n4999), .B0(n6532), .Y(n3383) );
  OAI2BB1X1 U7558 ( .A0N(N6429), .A1N(n4992), .B0(n6424), .Y(n3273) );
  OAI2BB1X1 U7559 ( .A0N(N5816), .A1N(n4990), .B0(n6078), .Y(n3660) );
  BUFX2 U7560 ( .A(reg_invalid2[1]), .Y(n5376) );
  INVX2 U7561 ( .A(reg_invalid2[4]), .Y(n7330) );
  INVX2 U7562 ( .A(reg_invalid2[0]), .Y(n7038) );
  OAI2BB1X1 U7563 ( .A0N(N5734), .A1N(n4989), .B0(n6174), .Y(n3770) );
  NAND2X1 U7564 ( .A(N5008), .B(n7177), .Y(n2665) );
  BUFX2 U7565 ( .A(reg_invalid2[3]), .Y(n5374) );
  OAI2BB1X1 U7566 ( .A0N(N5817), .A1N(n4990), .B0(n6077), .Y(n3659) );
  OR2X1 U7567 ( .A(reg_invalid2[0]), .B(n7035), .Y(n2804) );
  NAND2X1 U7568 ( .A(N5010), .B(n7177), .Y(n2664) );
  NAND3X1 U7569 ( .A(n5375), .B(n2715), .C(reg_invalid2[4]), .Y(n2705) );
  OAI2BB1X1 U7570 ( .A0N(N5775), .A1N(n4991), .B0(n6126), .Y(n3715) );
  OAI2BB1X1 U7571 ( .A0N(N5513), .A1N(n5002), .B0(n6272), .Y(n3879) );
  OAI2BB1X1 U7572 ( .A0N(N5776), .A1N(n4991), .B0(n6125), .Y(n3714) );
  OAI2BB1X1 U7573 ( .A0N(N5472), .A1N(n5003), .B0(n6323), .Y(n3925) );
  OAI2BB1X1 U7574 ( .A0N(N5431), .A1N(n5005), .B0(n5936), .Y(n3965) );
  OAI2BB1X1 U7575 ( .A0N(N5512), .A1N(n5002), .B0(n6273), .Y(n3880) );
  OR2X1 U7576 ( .A(reg_invalid2[0]), .B(n5376), .Y(n1910) );
  BUFX2 U7577 ( .A(reg_invalid2[5]), .Y(n5373) );
  INVX2 U7578 ( .A(n1434), .Y(n6390) );
  NOR4BX1 U7579 ( .AN(n2812), .B(reg_invalid2[7]), .C(reg_invalid2[8]), .D(
        n5373), .Y(n1434) );
  NOR3X1 U7580 ( .A(n7331), .B(reg_invalid2[4]), .C(n5374), .Y(n2812) );
  OAI2BB1X1 U7581 ( .A0N(N5430), .A1N(n5005), .B0(n5937), .Y(n3966) );
  OAI2BB1X1 U7582 ( .A0N(N5694), .A1N(n4998), .B0(n6222), .Y(n3824) );
  NAND2X1 U7583 ( .A(N5012), .B(n7177), .Y(n2659) );
  BUFX2 U7584 ( .A(reg_invalid2[2]), .Y(n5375) );
  OAI2BB1X1 U7585 ( .A0N(N6220), .A1N(n4995), .B0(n6703), .Y(n3552) );
  OAI2BB1X1 U7586 ( .A0N(N5471), .A1N(n5003), .B0(n6324), .Y(n3926) );
  OAI2BB1X1 U7587 ( .A0N(N5693), .A1N(n4998), .B0(n6223), .Y(n3825) );
  NAND2X1 U7588 ( .A(N5014), .B(n7177), .Y(n2658) );
  OAI2BB1X1 U7589 ( .A0N(N5815), .A1N(n4990), .B0(n6079), .Y(n3661) );
  OAI2BB1X1 U7590 ( .A0N(N6426), .A1N(n4992), .B0(n6427), .Y(n3276) );
  OAI2BB1X1 U7591 ( .A0N(N6221), .A1N(n4995), .B0(n6702), .Y(n3551) );
  INVX2 U7592 ( .A(reg_invalid2[6]), .Y(n7331) );
  OAI2BB1X1 U7593 ( .A0N(N6384), .A1N(n5000), .B0(n6482), .Y(n3332) );
  OAI2BB1X1 U7594 ( .A0N(N5733), .A1N(n4989), .B0(n6175), .Y(n3771) );
  OAI2BB1X1 U7595 ( .A0N(N6180), .A1N(n4994), .B0(n6757), .Y(n3606) );
  OAI2BB1X1 U7596 ( .A0N(N6385), .A1N(n5000), .B0(n6481), .Y(n3331) );
  OAI2BB1X1 U7597 ( .A0N(N6262), .A1N(n4996), .B0(n6647), .Y(n3496) );
  OAI2BB1X1 U7598 ( .A0N(N6303), .A1N(n4997), .B0(n6591), .Y(n3441) );
  OAI2BB1X1 U7599 ( .A0N(N5511), .A1N(n5002), .B0(n6274), .Y(n3881) );
  OAI2BB1X1 U7600 ( .A0N(N5774), .A1N(n4991), .B0(n6127), .Y(n3716) );
  OAI2BB1X1 U7601 ( .A0N(N6261), .A1N(n4996), .B0(n6648), .Y(n3497) );
  OAI2BB1X1 U7602 ( .A0N(N5470), .A1N(n5003), .B0(n6325), .Y(n3927) );
  OAI2BB1X1 U7603 ( .A0N(N5429), .A1N(n5005), .B0(n5938), .Y(n3967) );
  OAI2BB1X1 U7604 ( .A0N(N5732), .A1N(n4989), .B0(n6176), .Y(n3772) );
  OAI2BB1X1 U7605 ( .A0N(N5773), .A1N(n4991), .B0(n6128), .Y(n3717) );
  OAI2BB1X1 U7606 ( .A0N(N6302), .A1N(n4997), .B0(n6592), .Y(n3442) );
  OAI2BB1X1 U7607 ( .A0N(N6179), .A1N(n4994), .B0(n6758), .Y(n3607) );
  OAI2BB1X1 U7608 ( .A0N(N6344), .A1N(n4999), .B0(n6535), .Y(n3386) );
  OAI2BB1X1 U7609 ( .A0N(N6467), .A1N(n4993), .B0(n6373), .Y(n3221) );
  OAI2BB1X1 U7610 ( .A0N(N6425), .A1N(n4992), .B0(n6428), .Y(n3277) );
  OAI2BB1X1 U7611 ( .A0N(N6343), .A1N(n4999), .B0(n6536), .Y(n3387) );
  OAI2BB1X1 U7612 ( .A0N(N6466), .A1N(n4993), .B0(n6374), .Y(n3222) );
  OAI2BB1X1 U7613 ( .A0N(N5692), .A1N(n4998), .B0(n6224), .Y(n3826) );
  OAI2BB1X1 U7614 ( .A0N(N5510), .A1N(n5002), .B0(n6275), .Y(n3882) );
  OAI2BB1X1 U7615 ( .A0N(N5428), .A1N(n5005), .B0(n5939), .Y(n3968) );
  OAI2BB1X1 U7616 ( .A0N(N5469), .A1N(n5003), .B0(n6326), .Y(n3928) );
  OAI221X1 U7617 ( .A0(n7312), .A1(n2735), .B0(n7236), .B1(n2686), .C0(n2736), 
        .Y(N4784) );
  AOI222XL U7618 ( .A0(n2737), .A1(n5377), .B0(temp_i_mat_idx[3]), .B1(n2738), 
        .C0(n2739), .C1(count[13]), .Y(n2736) );
  NAND2X1 U7619 ( .A(in_valid), .B(n1314), .Y(n2539) );
  OAI2BB1X1 U7620 ( .A0N(N5814), .A1N(n4990), .B0(n6080), .Y(n3662) );
  NAND3X1 U7621 ( .A(n2769), .B(n2770), .C(n2771), .Y(N4779) );
  AOI221XL U7622 ( .A0(n2772), .A1(n7023), .B0(n7030), .B1(n2758), .C0(n2773), 
        .Y(n2771) );
  AOI22X1 U7623 ( .A0(n7190), .A1(N5059), .B0(n7233), .B1(i_mat_idx), .Y(n2769) );
  AOI222XL U7624 ( .A0(n2737), .A1(n5571), .B0(temp_i_mat_idx[0]), .B1(n2748), 
        .C0(n2739), .C1(N5061), .Y(n2770) );
  OAI2BB1X1 U7625 ( .A0N(N5691), .A1N(n4998), .B0(n6225), .Y(n3827) );
  OAI2BB1X1 U7626 ( .A0N(N5731), .A1N(n4989), .B0(n6177), .Y(n3773) );
  NAND2X1 U7627 ( .A(n2746), .B(n2747), .Y(N4782) );
  AOI221XL U7628 ( .A0(temp_i_mat_idx[3]), .A1(n2748), .B0(n2739), .B1(n5378), 
        .C0(n2749), .Y(n2747) );
  AOI222XL U7629 ( .A0(n7231), .A1(temp_i_mat_idx[0]), .B0(n2737), .B1(N5118), 
        .C0(n7190), .C1(n5568), .Y(n2746) );
  OAI22X1 U7630 ( .A0(n2750), .A1(n7236), .B0(n2744), .B1(n7235), .Y(n2749) );
  NAND2X1 U7631 ( .A(n2740), .B(n2741), .Y(N4783) );
  AOI222XL U7632 ( .A0(n2739), .A1(n5377), .B0(temp_i_mat_idx[2]), .B1(n7207), 
        .C0(temp_i_mat_idx[3]), .C1(n2743), .Y(n2741) );
  AOI222XL U7633 ( .A0(n7231), .A1(temp_i_mat_idx[1]), .B0(n2737), .B1(n5378), 
        .C0(n7190), .C1(N5118), .Y(n2740) );
  INVX2 U7634 ( .A(n2744), .Y(n7207) );
  NAND2X1 U7635 ( .A(n2751), .B(n2752), .Y(N4781) );
  AOI221XL U7636 ( .A0(temp_i_mat_idx[2]), .A1(n2748), .B0(n2739), .B1(N5118), 
        .C0(n2753), .Y(n2752) );
  AOI222XL U7637 ( .A0(n7231), .A1(i_mat_idx), .B0(n2737), .B1(n5568), .C0(
        n7190), .C1(N5061), .Y(n2751) );
  OAI22X1 U7638 ( .A0(n2750), .A1(n7235), .B0(n2744), .B1(n7234), .Y(n2753) );
  INVX2 U7639 ( .A(reg_matrix_size[3]), .Y(n7036) );
  OAI2BB1X1 U7640 ( .A0N(N5509), .A1N(n5002), .B0(n6276), .Y(n3883) );
  OAI2BB2X1 U7641 ( .B0(n1281), .B1(n7479), .A0N(N4935), .A1N(n7181), .Y(n3150) );
  OAI2BB2X1 U7642 ( .B0(n1281), .B1(n7475), .A0N(N4931), .A1N(n7181), .Y(n3154) );
  INVX2 U7643 ( .A(count58[2]), .Y(n7475) );
  OAI2BB2X1 U7644 ( .B0(n1281), .B1(n7474), .A0N(N4930), .A1N(n7181), .Y(n3155) );
  INVX2 U7645 ( .A(count58[1]), .Y(n7474) );
  OAI2BB2X1 U7646 ( .B0(n1281), .B1(n7473), .A0N(N4929), .A1N(n7181), .Y(n3156) );
  INVX2 U7647 ( .A(count58[0]), .Y(n7473) );
  OAI2BB2X1 U7648 ( .B0(n1224), .B1(n7444), .A0N(N4850), .A1N(n7184), .Y(n3115) );
  INVX2 U7649 ( .A(count08[6]), .Y(n7444) );
  OAI2BB2X1 U7650 ( .B0(n1224), .B1(n7443), .A0N(N4849), .A1N(n7184), .Y(n3116) );
  INVX2 U7651 ( .A(count08[5]), .Y(n7443) );
  OAI2BB2X1 U7652 ( .B0(n1224), .B1(n7442), .A0N(N4848), .A1N(n7184), .Y(n3117) );
  INVX2 U7653 ( .A(count08[4]), .Y(n7442) );
  OAI2BB2X1 U7654 ( .B0(n1224), .B1(n7441), .A0N(N4847), .A1N(n7184), .Y(n3118) );
  INVX2 U7655 ( .A(count08[3]), .Y(n7441) );
  OAI2BB2X1 U7656 ( .B0(n1224), .B1(n7440), .A0N(N4846), .A1N(n7184), .Y(n3119) );
  INVX2 U7657 ( .A(count08[2]), .Y(n7440) );
  OAI2BB2X1 U7658 ( .B0(n1224), .B1(n7439), .A0N(N4845), .A1N(n7184), .Y(n3120) );
  INVX2 U7659 ( .A(count08[1]), .Y(n7439) );
  OAI2BB2X1 U7660 ( .B0(n1224), .B1(n7438), .A0N(N4844), .A1N(n7184), .Y(n3121) );
  OAI2BB2X1 U7661 ( .B0(n1271), .B1(n7472), .A0N(N4918), .A1N(n7182), .Y(n3143) );
  OAI2BB2X1 U7662 ( .B0(n1271), .B1(n7468), .A0N(N4914), .A1N(n7182), .Y(n3147) );
  INVX2 U7663 ( .A(count48[2]), .Y(n7468) );
  OAI2BB2X1 U7664 ( .B0(n1271), .B1(n7467), .A0N(N4913), .A1N(n7182), .Y(n3148) );
  INVX2 U7665 ( .A(count48[1]), .Y(n7467) );
  OAI2BB2X1 U7666 ( .B0(n1271), .B1(n7466), .A0N(N4912), .A1N(n7182), .Y(n3149) );
  INVX2 U7667 ( .A(count48[0]), .Y(n7466) );
  OAI2BB2X1 U7668 ( .B0(n1238), .B1(n7451), .A0N(N4867), .A1N(n7183), .Y(n3122) );
  INVX2 U7669 ( .A(count18[6]), .Y(n7451) );
  OAI2BB2X1 U7670 ( .B0(n1238), .B1(n7450), .A0N(N4866), .A1N(n7183), .Y(n3123) );
  INVX2 U7671 ( .A(count18[5]), .Y(n7450) );
  OAI2BB2X1 U7672 ( .B0(n1238), .B1(n7449), .A0N(N4865), .A1N(n7183), .Y(n3124) );
  INVX2 U7673 ( .A(count18[4]), .Y(n7449) );
  OAI2BB2X1 U7674 ( .B0(n1238), .B1(n7448), .A0N(N4864), .A1N(n7183), .Y(n3125) );
  INVX2 U7675 ( .A(count18[3]), .Y(n7448) );
  OAI2BB2X1 U7676 ( .B0(n1238), .B1(n7447), .A0N(N4863), .A1N(n7183), .Y(n3126) );
  INVX2 U7677 ( .A(count18[2]), .Y(n7447) );
  OAI2BB2X1 U7678 ( .B0(n1238), .B1(n7446), .A0N(N4862), .A1N(n7183), .Y(n3127) );
  INVX2 U7679 ( .A(count18[1]), .Y(n7446) );
  OAI2BB2X1 U7680 ( .B0(n1238), .B1(n7445), .A0N(N4861), .A1N(n7183), .Y(n3128) );
  NAND2X1 U7681 ( .A(n2759), .B(n2760), .Y(N4780) );
  AOI221XL U7682 ( .A0(n2737), .A1(N5061), .B0(n7190), .B1(n5571), .C0(n2767), 
        .Y(n2759) );
  AOI221XL U7683 ( .A0(temp_i_mat_idx[1]), .A1(n2748), .B0(n2739), .B1(n5568), 
        .C0(n2761), .Y(n2760) );
  OAI2BB1X1 U7684 ( .A0N(i_mat_idx), .A1N(n7208), .B0(n2768), .Y(n2767) );
  OAI2BB2X1 U7685 ( .B0(n1248), .B1(n7458), .A0N(N4884), .A1N(n7180), .Y(n3129) );
  INVX2 U7686 ( .A(count28[6]), .Y(n7458) );
  OAI2BB2X1 U7687 ( .B0(n1248), .B1(n7457), .A0N(N4883), .A1N(n7180), .Y(n3130) );
  INVX2 U7688 ( .A(count28[5]), .Y(n7457) );
  OAI2BB2X1 U7689 ( .B0(n1248), .B1(n7456), .A0N(N4882), .A1N(n7180), .Y(n3131) );
  INVX2 U7690 ( .A(count28[4]), .Y(n7456) );
  OAI2BB2X1 U7691 ( .B0(n1248), .B1(n7455), .A0N(N4881), .A1N(n7180), .Y(n3132) );
  INVX2 U7692 ( .A(count28[3]), .Y(n7455) );
  OAI2BB2X1 U7693 ( .B0(n1248), .B1(n7454), .A0N(N4880), .A1N(n7180), .Y(n3133) );
  INVX2 U7694 ( .A(count28[2]), .Y(n7454) );
  OAI2BB2X1 U7695 ( .B0(n1248), .B1(n7453), .A0N(N4879), .A1N(n7180), .Y(n3134) );
  INVX2 U7696 ( .A(count28[1]), .Y(n7453) );
  OAI2BB2X1 U7697 ( .B0(n1248), .B1(n7452), .A0N(N4878), .A1N(n7180), .Y(n3135) );
  INVX2 U7698 ( .A(count28[0]), .Y(n7452) );
  OAI2BB2X1 U7699 ( .B0(n1292), .B1(n7486), .A0N(N4952), .A1N(n7179), .Y(n3157) );
  INVX2 U7700 ( .A(count68[6]), .Y(n7486) );
  OAI2BB2X1 U7701 ( .B0(n1292), .B1(n7485), .A0N(N4951), .A1N(n7179), .Y(n3158) );
  INVX2 U7702 ( .A(count68[5]), .Y(n7485) );
  OAI2BB2X1 U7703 ( .B0(n1292), .B1(n7484), .A0N(N4950), .A1N(n7179), .Y(n3159) );
  INVX2 U7704 ( .A(count68[4]), .Y(n7484) );
  OAI2BB2X1 U7705 ( .B0(n1292), .B1(n7483), .A0N(N4949), .A1N(n7179), .Y(n3160) );
  INVX2 U7706 ( .A(count68[3]), .Y(n7483) );
  OAI2BB2X1 U7707 ( .B0(n1292), .B1(n7482), .A0N(N4948), .A1N(n7179), .Y(n3161) );
  INVX2 U7708 ( .A(count68[2]), .Y(n7482) );
  OAI2BB2X1 U7709 ( .B0(n1292), .B1(n7481), .A0N(N4947), .A1N(n7179), .Y(n3162) );
  INVX2 U7710 ( .A(count68[1]), .Y(n7481) );
  OAI2BB2X1 U7711 ( .B0(n1292), .B1(n7480), .A0N(N4946), .A1N(n7179), .Y(n3163) );
  INVX2 U7712 ( .A(count68[0]), .Y(n7480) );
  INVX2 U7713 ( .A(reg_matrix_size[2]), .Y(n5574) );
  OAI2BB1X1 U7714 ( .A0N(N5427), .A1N(n5005), .B0(n5940), .Y(n3969) );
  OAI2BB1X1 U7715 ( .A0N(N5729), .A1N(n4989), .B0(n6179), .Y(n3775) );
  OAI2BB1X1 U7716 ( .A0N(N5468), .A1N(n5003), .B0(n6327), .Y(n3929) );
  OAI2BB1X1 U7717 ( .A0N(N5730), .A1N(n4989), .B0(n6178), .Y(n3774) );
  OAI2BB1X1 U7718 ( .A0N(N6258), .A1N(n4996), .B0(n6652), .Y(n3500) );
  OR2X1 U7719 ( .A(n6651), .B(n6661), .Y(n6652) );
  INVX2 U7720 ( .A(y_out_sum9[5]), .Y(n6651) );
  OAI2BB1X1 U7721 ( .A0N(N6217), .A1N(n4995), .B0(n6707), .Y(n3555) );
  OR2X1 U7722 ( .A(n6706), .B(n6716), .Y(n6707) );
  INVX2 U7723 ( .A(y_out_sum8[5]), .Y(n6706) );
  OAI2BB1X1 U7724 ( .A0N(N5813), .A1N(n4990), .B0(n6081), .Y(n3663) );
  OAI2BB1X1 U7725 ( .A0N(N5772), .A1N(n4991), .B0(n6129), .Y(n3718) );
  OAI2BB1X1 U7726 ( .A0N(N5690), .A1N(n4998), .B0(n6226), .Y(n3828) );
  OAI2BB1X1 U7727 ( .A0N(N5771), .A1N(n4991), .B0(n6130), .Y(n3719) );
  OAI2BB1X1 U7728 ( .A0N(N5812), .A1N(n4990), .B0(n6082), .Y(n3664) );
  OAI2BB1X1 U7729 ( .A0N(N5426), .A1N(n5005), .B0(n5941), .Y(n3970) );
  OAI2BB1X1 U7730 ( .A0N(N5508), .A1N(n5002), .B0(n6277), .Y(n3884) );
  OAI2BB1X1 U7731 ( .A0N(N5507), .A1N(n5002), .B0(n6278), .Y(n3885) );
  OAI2BB1X1 U7732 ( .A0N(N6176), .A1N(n4994), .B0(n6762), .Y(n3610) );
  OR2X1 U7733 ( .A(n6761), .B(n6771), .Y(n6762) );
  INVX2 U7734 ( .A(y_out_sum7[5]), .Y(n6761) );
  OAI2BB1X1 U7735 ( .A0N(N5467), .A1N(n5003), .B0(n6328), .Y(n3930) );
  OAI2BB1X1 U7736 ( .A0N(N6381), .A1N(n5000), .B0(n6486), .Y(n3335) );
  OR2X1 U7737 ( .A(n6485), .B(n6495), .Y(n6486) );
  INVX2 U7738 ( .A(y_out_sum12[5]), .Y(n6485) );
  OAI2BB2X1 U7739 ( .B0(n1302), .B1(n7493), .A0N(N4969), .A1N(n7178), .Y(n3164) );
  INVX2 U7740 ( .A(count78[6]), .Y(n7493) );
  OAI2BB2X1 U7741 ( .B0(n1302), .B1(n7492), .A0N(N4968), .A1N(n7178), .Y(n3165) );
  INVX2 U7742 ( .A(count78[5]), .Y(n7492) );
  OAI2BB2X1 U7743 ( .B0(n1302), .B1(n7491), .A0N(N4967), .A1N(n7178), .Y(n3166) );
  INVX2 U7744 ( .A(count78[4]), .Y(n7491) );
  OAI2BB2X1 U7745 ( .B0(n1302), .B1(n7490), .A0N(N4966), .A1N(n7178), .Y(n3167) );
  INVX2 U7746 ( .A(count78[3]), .Y(n7490) );
  OAI2BB2X1 U7747 ( .B0(n1302), .B1(n7489), .A0N(N4965), .A1N(n7178), .Y(n3168) );
  INVX2 U7748 ( .A(count78[2]), .Y(n7489) );
  OAI2BB2X1 U7749 ( .B0(n1302), .B1(n7488), .A0N(N4964), .A1N(n7178), .Y(n3169) );
  INVX2 U7750 ( .A(count78[1]), .Y(n7488) );
  OAI2BB2X1 U7751 ( .B0(n1302), .B1(n7487), .A0N(N4963), .A1N(n7178), .Y(n3170) );
  INVX2 U7752 ( .A(count78[0]), .Y(n7487) );
  OAI2BB2X1 U7753 ( .B0(n1259), .B1(n7465), .A0N(N4901), .A1N(n7185), .Y(n3136) );
  OAI2BB2X1 U7754 ( .B0(n1259), .B1(n7461), .A0N(N4897), .A1N(n7185), .Y(n3140) );
  INVX2 U7755 ( .A(count38[2]), .Y(n7461) );
  OAI2BB2X1 U7756 ( .B0(n1259), .B1(n7460), .A0N(N4896), .A1N(n7185), .Y(n3141) );
  INVX2 U7757 ( .A(count38[1]), .Y(n7460) );
  OAI2BB2X1 U7758 ( .B0(n1259), .B1(n7459), .A0N(N4895), .A1N(n7185), .Y(n3142) );
  INVX2 U7759 ( .A(count38[0]), .Y(n7459) );
  OAI2BB1X1 U7760 ( .A0N(N5689), .A1N(n4998), .B0(n6227), .Y(n3829) );
  OAI2BB1X1 U7761 ( .A0N(N6257), .A1N(n4996), .B0(n6654), .Y(n3501) );
  OR2X1 U7762 ( .A(n6653), .B(n6661), .Y(n6654) );
  INVX2 U7763 ( .A(y_out_sum9[4]), .Y(n6653) );
  OAI2BB1X1 U7764 ( .A0N(N6216), .A1N(n4995), .B0(n6709), .Y(n3556) );
  OR2X1 U7765 ( .A(n6708), .B(n6716), .Y(n6709) );
  INVX2 U7766 ( .A(y_out_sum8[4]), .Y(n6708) );
  OAI2BB2X1 U7767 ( .B0(n7303), .B1(n4848), .A0N(N4584), .A1N(n2376), .Y(n4025) );
  OAI2BB2X1 U7768 ( .B0(n7315), .B1(n4848), .A0N(N4599), .A1N(n2376), .Y(n4011) );
  OAI2BB2X1 U7769 ( .B0(n7314), .B1(n4848), .A0N(N4598), .A1N(n2376), .Y(n4012) );
  INVX2 U7770 ( .A(count[14]), .Y(n7314) );
  INVX2 U7771 ( .A(in_valid), .Y(n7168) );
  NOR3X1 U7772 ( .A(reg_matrix_size[2]), .B(reg_matrix_size[3]), .C(n7037), 
        .Y(n117) );
  OAI2BB1X1 U7773 ( .A0N(N5688), .A1N(n4998), .B0(n6228), .Y(n3830) );
  INVX2 U7774 ( .A(reg_matrix_size[1]), .Y(n7037) );
  OAI2BB1X1 U7775 ( .A0N(N6422), .A1N(n4992), .B0(n6432), .Y(n3280) );
  OR2X1 U7776 ( .A(n6431), .B(n6441), .Y(n6432) );
  INVX2 U7777 ( .A(y_out_sum13[5]), .Y(n6431) );
  AND2X1 U7778 ( .A(D1[119]), .B(n5422), .Y(N5378) );
  AND2X1 U7779 ( .A(D1[118]), .B(n5422), .Y(N5377) );
  AND2X1 U7780 ( .A(D1[117]), .B(n5422), .Y(N5376) );
  AND2X1 U7781 ( .A(D1[116]), .B(n5422), .Y(N5375) );
  AND2X1 U7782 ( .A(D1[115]), .B(n5422), .Y(N5374) );
  AND2X1 U7783 ( .A(D1[114]), .B(n5422), .Y(N5373) );
  AND2X1 U7784 ( .A(D1[113]), .B(n5422), .Y(N5372) );
  AND2X1 U7785 ( .A(D1[112]), .B(n5422), .Y(N5371) );
  AND2X1 U7786 ( .A(D1[111]), .B(n5422), .Y(N5370) );
  AND2X1 U7787 ( .A(D1[110]), .B(n5422), .Y(N5369) );
  AND2X1 U7788 ( .A(D1[109]), .B(n5422), .Y(N5368) );
  AND2X1 U7789 ( .A(D1[108]), .B(n5422), .Y(N5367) );
  AND2X1 U7790 ( .A(D1[107]), .B(n5422), .Y(N5366) );
  AND2X1 U7791 ( .A(D1[106]), .B(n5422), .Y(N5365) );
  AND2X1 U7792 ( .A(D1[105]), .B(n5422), .Y(N5364) );
  AND2X1 U7793 ( .A(D1[104]), .B(n5422), .Y(N5363) );
  AND2X1 U7794 ( .A(D1[103]), .B(n5422), .Y(N5362) );
  AND2X1 U7795 ( .A(D1[102]), .B(n5422), .Y(N5361) );
  AND2X1 U7796 ( .A(D1[101]), .B(n5422), .Y(N5360) );
  AND2X1 U7797 ( .A(D1[100]), .B(n5418), .Y(N5359) );
  AND2X1 U7798 ( .A(D1[99]), .B(n5416), .Y(N5358) );
  AND2X1 U7799 ( .A(D1[98]), .B(n5422), .Y(N5357) );
  AND2X1 U7800 ( .A(D1[97]), .B(n5418), .Y(N5356) );
  AND2X1 U7801 ( .A(D1[96]), .B(n5416), .Y(N5355) );
  AND2X1 U7802 ( .A(D1[95]), .B(n5421), .Y(N5354) );
  AND2X1 U7803 ( .A(D1[94]), .B(n5421), .Y(N5353) );
  AND2X1 U7804 ( .A(D1[93]), .B(n5421), .Y(N5352) );
  AND2X1 U7805 ( .A(D1[92]), .B(n5421), .Y(N5351) );
  AND2X1 U7806 ( .A(D1[91]), .B(n5421), .Y(N5350) );
  AND2X1 U7807 ( .A(D1[90]), .B(n5421), .Y(N5349) );
  AND2X1 U7808 ( .A(D1[89]), .B(n5421), .Y(N5348) );
  AND2X1 U7809 ( .A(D1[88]), .B(n5421), .Y(N5347) );
  AND2X1 U7810 ( .A(D1[87]), .B(n5421), .Y(N5346) );
  AND2X1 U7811 ( .A(D1[86]), .B(n5421), .Y(N5345) );
  AND2X1 U7812 ( .A(D1[85]), .B(n5421), .Y(N5344) );
  AND2X1 U7813 ( .A(D1[84]), .B(n5421), .Y(N5343) );
  AND2X1 U7814 ( .A(D1[83]), .B(n5420), .Y(N5342) );
  AND2X1 U7815 ( .A(D1[82]), .B(n5420), .Y(N5341) );
  AND2X1 U7816 ( .A(D1[81]), .B(n5420), .Y(N5340) );
  AND2X1 U7817 ( .A(D1[80]), .B(n5420), .Y(N5339) );
  AND2X1 U7818 ( .A(D1[79]), .B(n5420), .Y(N5338) );
  AND2X1 U7819 ( .A(D1[78]), .B(n5420), .Y(N5337) );
  AND2X1 U7820 ( .A(D1[77]), .B(n5420), .Y(N5336) );
  AND2X1 U7821 ( .A(D1[76]), .B(n5420), .Y(N5335) );
  AND2X1 U7822 ( .A(D1[75]), .B(n5420), .Y(N5334) );
  AND2X1 U7823 ( .A(D1[74]), .B(n5420), .Y(N5333) );
  AND2X1 U7824 ( .A(D1[73]), .B(n5420), .Y(N5332) );
  AND2X1 U7825 ( .A(D1[72]), .B(n5420), .Y(N5331) );
  AND2X1 U7826 ( .A(D1[71]), .B(n5419), .Y(N5330) );
  AND2X1 U7827 ( .A(D1[70]), .B(n5419), .Y(N5329) );
  AND2X1 U7828 ( .A(D1[69]), .B(n5419), .Y(N5328) );
  AND2X1 U7829 ( .A(D1[68]), .B(n5419), .Y(N5327) );
  AND2X1 U7830 ( .A(D1[67]), .B(n5419), .Y(N5326) );
  AND2X1 U7831 ( .A(D1[66]), .B(n5419), .Y(N5325) );
  AND2X1 U7832 ( .A(D1[65]), .B(n5419), .Y(N5324) );
  AND2X1 U7833 ( .A(D1[64]), .B(n5419), .Y(N5323) );
  AND2X1 U7834 ( .A(D1[63]), .B(n5419), .Y(N5322) );
  AND2X1 U7835 ( .A(D1[62]), .B(n5419), .Y(N5321) );
  AND2X1 U7836 ( .A(D1[61]), .B(n5419), .Y(N5320) );
  AND2X1 U7837 ( .A(D1[60]), .B(n5419), .Y(N5319) );
  AND2X1 U7838 ( .A(D1[59]), .B(n5418), .Y(N5318) );
  AND2X1 U7839 ( .A(D1[58]), .B(n5418), .Y(N5317) );
  AND2X1 U7840 ( .A(D1[57]), .B(n5418), .Y(N5316) );
  AND2X1 U7841 ( .A(D1[56]), .B(n5418), .Y(N5315) );
  AND2X1 U7842 ( .A(D1[55]), .B(n5418), .Y(N5314) );
  AND2X1 U7843 ( .A(D1[54]), .B(n5418), .Y(N5313) );
  AND2X1 U7844 ( .A(D1[53]), .B(n5418), .Y(N5312) );
  AND2X1 U7845 ( .A(D1[52]), .B(n5418), .Y(N5311) );
  AND2X1 U7846 ( .A(D1[51]), .B(n5418), .Y(N5310) );
  AND2X1 U7847 ( .A(D1[50]), .B(n5418), .Y(N5309) );
  AND2X1 U7848 ( .A(D1[49]), .B(n5418), .Y(N5308) );
  AND2X1 U7849 ( .A(D1[48]), .B(n5418), .Y(N5307) );
  AND2X1 U7850 ( .A(D1[47]), .B(n5418), .Y(N5306) );
  AND2X1 U7851 ( .A(D1[46]), .B(n5418), .Y(N5305) );
  AND2X1 U7852 ( .A(D1[45]), .B(n5418), .Y(N5304) );
  AND2X1 U7853 ( .A(D1[44]), .B(n5418), .Y(N5303) );
  AND2X1 U7854 ( .A(D1[43]), .B(n5418), .Y(N5302) );
  AND2X1 U7855 ( .A(D1[42]), .B(n5418), .Y(N5301) );
  AND2X1 U7856 ( .A(D1[41]), .B(n5418), .Y(N5300) );
  AND2X1 U7857 ( .A(D1[40]), .B(n5418), .Y(N5299) );
  AND2X1 U7858 ( .A(D1[39]), .B(n5418), .Y(N5298) );
  AND2X1 U7859 ( .A(D1[38]), .B(n5418), .Y(N5297) );
  AND2X1 U7860 ( .A(D1[37]), .B(n5418), .Y(N5296) );
  AND2X1 U7861 ( .A(D1[36]), .B(n5418), .Y(N5295) );
  AND2X1 U7862 ( .A(D1[35]), .B(n5417), .Y(N5294) );
  AND2X1 U7863 ( .A(D1[34]), .B(n5417), .Y(N5293) );
  AND2X1 U7864 ( .A(D1[33]), .B(n5417), .Y(N5292) );
  AND2X1 U7865 ( .A(D1[32]), .B(n5417), .Y(N5291) );
  AND2X1 U7866 ( .A(D1[31]), .B(n5417), .Y(N5290) );
  AND2X1 U7867 ( .A(D1[30]), .B(n5417), .Y(N5289) );
  AND2X1 U7868 ( .A(D1[29]), .B(n5417), .Y(N5288) );
  AND2X1 U7869 ( .A(D1[28]), .B(n5417), .Y(N5287) );
  AND2X1 U7870 ( .A(D1[27]), .B(n5417), .Y(N5286) );
  AND2X1 U7871 ( .A(D1[26]), .B(n5417), .Y(N5285) );
  AND2X1 U7872 ( .A(D1[25]), .B(n5417), .Y(N5284) );
  AND2X1 U7873 ( .A(D1[24]), .B(n5417), .Y(N5283) );
  AND2X1 U7874 ( .A(D1[23]), .B(n5418), .Y(N5282) );
  AND2X1 U7875 ( .A(D1[22]), .B(n5418), .Y(N5281) );
  AND2X1 U7876 ( .A(D1[21]), .B(n5417), .Y(N5280) );
  AND2X1 U7877 ( .A(D1[20]), .B(n5422), .Y(N5279) );
  AND2X1 U7878 ( .A(D1[19]), .B(n5418), .Y(N5278) );
  AND2X1 U7879 ( .A(D1[18]), .B(n5418), .Y(N5277) );
  AND2X1 U7880 ( .A(D1[17]), .B(n5417), .Y(N5276) );
  AND2X1 U7881 ( .A(D1[16]), .B(n5422), .Y(N5275) );
  AND2X1 U7882 ( .A(D1[15]), .B(n5418), .Y(N5274) );
  AND2X1 U7883 ( .A(D1[14]), .B(n5418), .Y(N5273) );
  AND2X1 U7884 ( .A(D1[13]), .B(n5417), .Y(N5272) );
  AND2X1 U7885 ( .A(D1[12]), .B(n5422), .Y(N5271) );
  AND2X1 U7886 ( .A(D1[11]), .B(n5416), .Y(N5270) );
  AND2X1 U7887 ( .A(D1[10]), .B(n5416), .Y(N5269) );
  AND2X1 U7888 ( .A(D1[9]), .B(n5416), .Y(N5268) );
  AND2X1 U7889 ( .A(D1[8]), .B(n5416), .Y(N5267) );
  AND2X1 U7890 ( .A(D1[7]), .B(n5416), .Y(N5266) );
  AND2X1 U7891 ( .A(D1[6]), .B(n5416), .Y(N5265) );
  AND2X1 U7892 ( .A(D1[5]), .B(n5416), .Y(N5264) );
  AND2X1 U7893 ( .A(D1[4]), .B(n5416), .Y(N5263) );
  AND2X1 U7894 ( .A(D1[3]), .B(n5416), .Y(N5262) );
  AND2X1 U7895 ( .A(D1[2]), .B(n5416), .Y(N5261) );
  AND2X1 U7896 ( .A(D1[1]), .B(n5416), .Y(N5260) );
  AND2X1 U7897 ( .A(D1[0]), .B(n5416), .Y(N5259) );
  OAI2BB1X1 U7898 ( .A0N(N5770), .A1N(n4991), .B0(n6131), .Y(n3720) );
  OAI2BB1X1 U7899 ( .A0N(N5811), .A1N(n4990), .B0(n6083), .Y(n3665) );
  OAI2BB1X1 U7900 ( .A0N(N6340), .A1N(n4999), .B0(n6540), .Y(n3390) );
  OR2X1 U7901 ( .A(n6539), .B(n6549), .Y(n6540) );
  INVX2 U7902 ( .A(y_out_sum11[5]), .Y(n6539) );
  OAI2BB1X1 U7903 ( .A0N(N6299), .A1N(n4997), .B0(n6596), .Y(n3445) );
  OR2X1 U7904 ( .A(n6595), .B(n6605), .Y(n6596) );
  INVX2 U7905 ( .A(y_out_sum10[5]), .Y(n6595) );
  OAI2BB1X1 U7906 ( .A0N(N6463), .A1N(n4993), .B0(n6378), .Y(n3225) );
  OR2X1 U7907 ( .A(n6377), .B(n6387), .Y(n6378) );
  INVX2 U7908 ( .A(y_out_sum14[5]), .Y(n6377) );
  OAI2BB1X1 U7909 ( .A0N(N5425), .A1N(n5005), .B0(n5942), .Y(n3971) );
  AND2X1 U7910 ( .A(D1[126]), .B(n5417), .Y(N5385) );
  AND2X1 U7911 ( .A(D1[125]), .B(n5416), .Y(N5384) );
  AND2X1 U7912 ( .A(D1[124]), .B(n5422), .Y(N5383) );
  AND2X1 U7913 ( .A(D1[123]), .B(n5422), .Y(N5382) );
  AND2X1 U7914 ( .A(D1[122]), .B(n5422), .Y(N5381) );
  AND2X1 U7915 ( .A(D1[121]), .B(n5416), .Y(N5380) );
  AND2X1 U7916 ( .A(D1[120]), .B(n5422), .Y(N5379) );
  INVX2 U7917 ( .A(in_valid2), .Y(n7191) );
  NAND2X1 U7918 ( .A(n7203), .B(n2363), .Y(n2362) );
  OAI2BB1X1 U7919 ( .A0N(n7316), .A1N(reg_invalid2_signal), .B0(n7191), .Y(
        n2363) );
  INVX2 U7920 ( .A(N4685), .Y(n7316) );
  OAI2BB1X1 U7921 ( .A0N(N5466), .A1N(n5003), .B0(n6329), .Y(n3931) );
  OAI2BB1X1 U7922 ( .A0N(N5728), .A1N(n4989), .B0(n6180), .Y(n3776) );
  OAI2BB2X1 U7923 ( .B0(n7038), .B1(n2354), .A0N(N4694), .A1N(n7042), .Y(n3999) );
  NAND2X1 U7924 ( .A(in_valid), .B(in_slut), .Y(n132) );
  INVX2 U7925 ( .A(n135), .Y(n7169) );
  AOI32X1 U7926 ( .A0(matrix_size[0]), .A1(n7193), .A2(n7170), .B0(n132), .B1(
        reg_matrix_size[2]), .Y(n135) );
  OAI2BB2X1 U7927 ( .B0(n2354), .B1(n7333), .A0N(N4702), .A1N(n7042), .Y(n3992) );
  INVX2 U7928 ( .A(reg_invalid2[8]), .Y(n7333) );
  OAI2BB2X1 U7929 ( .B0(n2354), .B1(n7332), .A0N(N4701), .A1N(n7042), .Y(n3993) );
  INVX2 U7930 ( .A(reg_invalid2[7]), .Y(n7332) );
  OAI2BB1X1 U7931 ( .A0N(N5810), .A1N(n4990), .B0(n6084), .Y(n3666) );
  NAND2X1 U7932 ( .A(current_state[0]), .B(current_state[1]), .Y(n96) );
  OAI2BB1X1 U7933 ( .A0N(N5505), .A1N(n5002), .B0(n6280), .Y(n3887) );
  OAI222X1 U7934 ( .A0(n177), .A1(n178), .B0(n179), .B1(n5363), .C0(n181), 
        .C1(n182), .Y(n166) );
  AOI22X1 U7935 ( .A0(n5364), .A1(n7249), .B0(reg_length10[1]), .B1(n7254), 
        .Y(n181) );
  AOI221XL U7936 ( .A0(reg_length12[2]), .A1(n7255), .B0(reg_length12[1]), 
        .B1(n7254), .C0(n187), .Y(n177) );
  AOI21X1 U7937 ( .A0(n7041), .A1(n185), .B0(n186), .Y(n179) );
  OAI2BB1X1 U7938 ( .A0N(N5727), .A1N(n4989), .B0(n6181), .Y(n3777) );
  OAI2BB1X1 U7939 ( .A0N(N6421), .A1N(n4992), .B0(n6434), .Y(n3281) );
  OR2X1 U7940 ( .A(n6433), .B(n6441), .Y(n6434) );
  INVX2 U7941 ( .A(y_out_sum13[4]), .Y(n6433) );
  OAI2BB1X1 U7942 ( .A0N(N5769), .A1N(n4991), .B0(n6132), .Y(n3721) );
  OAI2BB1X1 U7943 ( .A0N(N6298), .A1N(n4997), .B0(n6598), .Y(n3446) );
  OR2X1 U7944 ( .A(n6597), .B(n6605), .Y(n6598) );
  INVX2 U7945 ( .A(y_out_sum10[4]), .Y(n6597) );
  OAI2BB1X1 U7946 ( .A0N(N6175), .A1N(n4994), .B0(n6764), .Y(n3611) );
  OR2X1 U7947 ( .A(n6763), .B(n6771), .Y(n6764) );
  INVX2 U7948 ( .A(y_out_sum7[4]), .Y(n6763) );
  OAI2BB1X1 U7949 ( .A0N(N6380), .A1N(n5000), .B0(n6488), .Y(n3336) );
  OR2X1 U7950 ( .A(n6487), .B(n6495), .Y(n6488) );
  INVX2 U7951 ( .A(y_out_sum12[4]), .Y(n6487) );
  OAI2BB1X1 U7952 ( .A0N(N6339), .A1N(n4999), .B0(n6542), .Y(n3391) );
  OR2X1 U7953 ( .A(n6541), .B(n6549), .Y(n6542) );
  INVX2 U7954 ( .A(y_out_sum11[4]), .Y(n6541) );
  OAI2BB1X1 U7955 ( .A0N(N6462), .A1N(n4993), .B0(n6380), .Y(n3226) );
  OR2X1 U7956 ( .A(n6379), .B(n6387), .Y(n6380) );
  INVX2 U7957 ( .A(y_out_sum14[4]), .Y(n6379) );
  OAI2BB1X1 U7958 ( .A0N(N5687), .A1N(n4998), .B0(n6229), .Y(n3831) );
  OAI2BB1X1 U7959 ( .A0N(N5465), .A1N(n5003), .B0(n6330), .Y(n3932) );
  OAI2BB1X1 U7960 ( .A0N(N5424), .A1N(n5005), .B0(n5943), .Y(n3972) );
  OAI2BB1X1 U7961 ( .A0N(N5506), .A1N(n5002), .B0(n6279), .Y(n3886) );
  INVX2 U7962 ( .A(matrix_size[1]), .Y(n7193) );
  OAI32X1 U7963 ( .A0(n132), .A1(matrix_size[0]), .A2(matrix_size[1]), .B0(
        n7170), .B1(n7037), .Y(n2850) );
  OAI2BB1X1 U7964 ( .A0N(N5686), .A1N(n4998), .B0(n6230), .Y(n3832) );
  OAI2BB1X1 U7965 ( .A0N(N5809), .A1N(n4990), .B0(n6085), .Y(n3667) );
  NAND2X1 U7966 ( .A(N7980), .B(reg_length14[0]), .Y(n297) );
  AOI222XL U7967 ( .A0(reg_length14[0]), .A1(n7248), .B0(n279), .B1(n280), 
        .C0(n7279), .C1(n282), .Y(n277) );
  OAI222X1 U7968 ( .A0(n283), .A1(n7594), .B0(n190), .B1(n7595), .C0(n188), 
        .C1(n7593), .Y(n282) );
  INVX2 U7969 ( .A(n343), .Y(n7248) );
  OAI222X1 U7970 ( .A0(n287), .A1(n7536), .B0(N7983), .B1(n289), .C0(n290), 
        .C1(n5016), .Y(n280) );
  AOI221XL U7971 ( .A0(y_out_sum14[5]), .A1(n300), .B0(y_out_sum14[4]), .B1(
        n301), .C0(n321), .Y(n6949) );
  OAI22X1 U7972 ( .A0(n297), .A1(n4907), .B0(n295), .B1(n4855), .Y(n321) );
  AOI32X1 U7973 ( .A0(n7535), .A1(n5016), .A2(n306), .B0(N7982), .B1(n307), 
        .Y(n289) );
  OAI22X1 U7974 ( .A0(n308), .A1(n7534), .B0(N7981), .B1(n309), .Y(n307) );
  OAI22X1 U7975 ( .A0(N7981), .A1(n6950), .B0(n7534), .B1(n6949), .Y(n306) );
  AOI221XL U7976 ( .A0(y_out_sum14[13]), .A1(n300), .B0(y_out_sum14[12]), .B1(
        n301), .C0(n313), .Y(n308) );
  AOI221XL U7977 ( .A0(y_out_sum14[1]), .A1(n300), .B0(y_out_sum14[0]), .B1(
        n301), .C0(n6948), .Y(n6950) );
  OAI22X1 U7978 ( .A0(n295), .A1(n4858), .B0(n297), .B1(n4906), .Y(n6948) );
  OAI2BB1X1 U7979 ( .A0N(N5423), .A1N(n5005), .B0(n5944), .Y(n3973) );
  OAI2BB1X1 U7980 ( .A0N(N5464), .A1N(n5003), .B0(n6331), .Y(n3933) );
  NOR3BX1 U7981 ( .AN(n2525), .B(next[3]), .C(n7292), .Y(n2531) );
  NOR4X1 U7982 ( .A(next[4]), .B(next[5]), .C(next[6]), .D(next[7]), .Y(n2525)
         );
  OAI211X1 U7983 ( .A0(n788), .A1(n7242), .B0(n790), .C0(n791), .Y(n787) );
  NOR4X1 U7984 ( .A(n809), .B(n5365), .C(reg_length12[2]), .D(reg_length12[1]), 
        .Y(n788) );
  INVX2 U7985 ( .A(n598), .Y(n7242) );
  AOI32X1 U7986 ( .A0(n802), .A1(n7047), .A2(n185), .B0(n211), .B1(n804), .Y(
        n790) );
  NOR3BX1 U7987 ( .AN(next[1]), .B(n5898), .C(n5897), .Y(n5015) );
  INVX2 U7988 ( .A(n5015), .Y(n171) );
  NAND3X1 U7989 ( .A(n929), .B(n7529), .C(shift[0]), .Y(n190) );
  NOR2X1 U7990 ( .A(shift[2]), .B(shift[3]), .Y(n923) );
  NOR2X1 U7991 ( .A(shift[4]), .B(shift[5]), .Y(n925) );
  AOI221XL U7992 ( .A0(y_out_sum14[9]), .A1(n300), .B0(y_out_sum14[8]), .B1(
        n301), .C0(n310), .Y(n309) );
  OAI22X1 U7993 ( .A0(n297), .A1(n4911), .B0(n295), .B1(n4860), .Y(n310) );
  NAND4X1 U7994 ( .A(shift[2]), .B(n7258), .C(n925), .D(n7531), .Y(n188) );
  INVX2 U7995 ( .A(shift[1]), .Y(n7529) );
  OAI22X1 U7996 ( .A0(n828), .A1(n5363), .B0(n829), .B1(n7241), .Y(n827) );
  NOR4X1 U7997 ( .A(n832), .B(reg_length14[0]), .C(reg_length14[2]), .D(
        reg_length14[1]), .Y(n829) );
  AOI221XL U7998 ( .A0(n185), .A1(n835), .B0(n7264), .B1(n836), .C0(n837), .Y(
        n828) );
  INVX2 U7999 ( .A(n279), .Y(n7241) );
  INVX2 U8000 ( .A(shift[0]), .Y(n7259) );
  NAND3X1 U8001 ( .A(n929), .B(n7259), .C(shift[1]), .Y(n283) );
  OAI2BB2X1 U8002 ( .B0(n7191), .B1(n7239), .A0N(n7191), .A1N(
        temp_w_mat_idx[3]), .Y(n2842) );
  OAI2BB2X1 U8003 ( .B0(n7191), .B1(n7236), .A0N(n7191), .A1N(
        temp_i_mat_idx[3]), .Y(n2846) );
  OAI2BB1X1 U8004 ( .A0N(N5768), .A1N(n4991), .B0(n6133), .Y(n3722) );
  OAI2BB1X1 U8005 ( .A0N(N5504), .A1N(n5002), .B0(n6282), .Y(n3888) );
  OR2X1 U8006 ( .A(n6286), .B(n6281), .Y(n6282) );
  INVX2 U8007 ( .A(y_out_sum2[2]), .Y(n6281) );
  INVX2 U8008 ( .A(next[2]), .Y(n7292) );
  AOI222XL U8009 ( .A0(n197), .A1(n198), .B0(n199), .B1(n200), .C0(n7272), 
        .C1(n202), .Y(n196) );
  OAI221X1 U8010 ( .A0(n5361), .A1(n7583), .B0(n5362), .B1(n7582), .C0(n210), 
        .Y(n200) );
  OAI221X1 U8011 ( .A0(n5361), .A1(n7564), .B0(n5362), .B1(n7563), .C0(n207), 
        .Y(n202) );
  AOI222XL U8012 ( .A0(reg_length9[3]), .A1(n7257), .B0(reg_length9[5]), .B1(
        n7260), .C0(reg_length9[4]), .C1(n7244), .Y(n210) );
  OAI22X1 U8013 ( .A0(n7191), .A1(n7234), .B0(in_valid2), .B1(n7235), .Y(n2848) );
  OAI22X1 U8014 ( .A0(n7191), .A1(n7235), .B0(in_valid2), .B1(n7236), .Y(n2847) );
  OAI22X1 U8015 ( .A0(n7191), .A1(n7238), .B0(in_valid2), .B1(n7239), .Y(n2843) );
  OAI22X1 U8016 ( .A0(n7191), .A1(n7237), .B0(in_valid2), .B1(n7238), .Y(n2844) );
  AOI22X1 U8017 ( .A0(N7982), .A1(n324), .B0(n325), .B1(n7535), .Y(n287) );
  OAI22X1 U8018 ( .A0(n326), .A1(n7534), .B0(N7981), .B1(n327), .Y(n325) );
  OAI22X1 U8019 ( .A0(n334), .A1(n7534), .B0(N7981), .B1(n335), .Y(n324) );
  AOI221XL U8020 ( .A0(y_out_sum14[17]), .A1(n300), .B0(y_out_sum14[16]), .B1(
        n301), .C0(n328), .Y(n327) );
  AOI221XL U8021 ( .A0(y_out_sum14[26]), .A1(n6947), .B0(y_out_sum14[27]), 
        .B1(n6956), .C0(n6943), .Y(n335) );
  OAI22X1 U8022 ( .A0(n6960), .A1(n6942), .B0(n6958), .B1(n6941), .Y(n6943) );
  AOI221XL U8023 ( .A0(y_out_sum14[22]), .A1(n6947), .B0(y_out_sum14[23]), 
        .B1(n6956), .C0(n6946), .Y(n326) );
  OAI22X1 U8024 ( .A0(n6960), .A1(n6945), .B0(n6958), .B1(n6944), .Y(n6946) );
  NAND2X1 U8025 ( .A(N7872), .B(reg_length11[0]), .Y(n361) );
  AOI222XL U8026 ( .A0(n346), .A1(n347), .B0(reg_length13[1]), .B1(n7253), 
        .C0(n349), .C1(n350), .Y(n275) );
  INVX2 U8027 ( .A(n407), .Y(n7253) );
  OAI222X1 U8028 ( .A0(n408), .A1(n7590), .B0(N7767), .B1(n410), .C0(n411), 
        .C1(n5018), .Y(n347) );
  OAI222X1 U8029 ( .A0(n351), .A1(n7562), .B0(N7875), .B1(n353), .C0(n354), 
        .C1(n5020), .Y(n350) );
  AOI221XL U8030 ( .A0(y_out_sum11[5]), .A1(n364), .B0(y_out_sum11[4]), .B1(
        n365), .C0(n385), .Y(n6925) );
  OAI22X1 U8031 ( .A0(n361), .A1(n4904), .B0(n359), .B1(n4852), .Y(n385) );
  AOI32X1 U8032 ( .A0(n7561), .A1(n5020), .A2(n370), .B0(N7874), .B1(n371), 
        .Y(n353) );
  OAI22X1 U8033 ( .A0(n372), .A1(n7560), .B0(N7873), .B1(n373), .Y(n371) );
  OAI22X1 U8034 ( .A0(N7873), .A1(n6926), .B0(n7560), .B1(n6925), .Y(n370) );
  AOI221XL U8035 ( .A0(y_out_sum11[13]), .A1(n364), .B0(y_out_sum11[12]), .B1(
        n365), .C0(n377), .Y(n372) );
  AOI2BB1X1 U8036 ( .A0N(reg_invalid2_signal), .A1N(in_valid2), .B0(n2365), 
        .Y(n4001) );
  NAND2X1 U8037 ( .A(N7764), .B(reg_length8[0]), .Y(n418) );
  AOI221XL U8038 ( .A0(y_out_sum8[5]), .A1(n421), .B0(y_out_sum8[4]), .B1(n422), .C0(n442), .Y(n6901) );
  OAI22X1 U8039 ( .A0(n418), .A1(n4914), .B0(n416), .B1(n4862), .Y(n442) );
  AOI32X1 U8040 ( .A0(n7589), .A1(n5018), .A2(n427), .B0(N7766), .B1(n428), 
        .Y(n410) );
  OAI22X1 U8041 ( .A0(n429), .A1(n7588), .B0(N7765), .B1(n430), .Y(n428) );
  OAI22X1 U8042 ( .A0(N7765), .A1(n6902), .B0(n7588), .B1(n6901), .Y(n427) );
  AOI221XL U8043 ( .A0(y_out_sum8[13]), .A1(n421), .B0(y_out_sum8[12]), .B1(
        n422), .C0(n434), .Y(n429) );
  AOI221XL U8044 ( .A0(y_out_sum14[30]), .A1(n6947), .B0(y_out_sum14[31]), 
        .B1(n6956), .C0(n6940), .Y(n334) );
  OAI22X1 U8045 ( .A0(n6960), .A1(n6939), .B0(n6958), .B1(n6938), .Y(n6940) );
  AOI221XL U8046 ( .A0(y_out_sum11[1]), .A1(n364), .B0(y_out_sum11[0]), .B1(
        n365), .C0(n6924), .Y(n6926) );
  OAI22X1 U8047 ( .A0(n359), .A1(n4853), .B0(n361), .B1(n4903), .Y(n6924) );
  AOI221XL U8048 ( .A0(y_out_sum8[1]), .A1(n421), .B0(y_out_sum8[0]), .B1(n422), .C0(n6900), .Y(n6902) );
  OAI22X1 U8049 ( .A0(n416), .A1(n4863), .B0(n418), .B1(n4913), .Y(n6900) );
  OAI2BB2X1 U8050 ( .B0(in_valid2), .B1(n7237), .A0N(in_valid2), .A1N(
        w_mat_idx), .Y(n2845) );
  OAI2BB2X1 U8051 ( .B0(in_valid2), .B1(n7234), .A0N(in_valid2), .A1N(
        i_mat_idx), .Y(n2849) );
  NOR2X1 U8052 ( .A(reg_length14[0]), .B(N7980), .Y(n300) );
  OAI2BB1X1 U8053 ( .A0N(N5463), .A1N(n5003), .B0(n6332), .Y(n3934) );
  AND2X1 U8054 ( .A(D3[14]), .B(in_valid), .Y(N5402) );
  AND2X1 U8055 ( .A(D3[13]), .B(in_valid), .Y(N5401) );
  AND2X1 U8056 ( .A(D3[12]), .B(in_valid), .Y(N5400) );
  AND2X1 U8057 ( .A(D3[11]), .B(in_valid), .Y(N5399) );
  AND2X1 U8058 ( .A(D3[10]), .B(in_valid), .Y(N5398) );
  AND2X1 U8059 ( .A(D3[9]), .B(in_valid), .Y(N5397) );
  AND2X1 U8060 ( .A(D3[8]), .B(in_valid), .Y(N5396) );
  AND2X1 U8061 ( .A(D3[7]), .B(in_valid), .Y(N5395) );
  AND2X1 U8062 ( .A(D3[6]), .B(in_valid), .Y(N5394) );
  AND2X1 U8063 ( .A(D3[5]), .B(in_valid), .Y(N5393) );
  AND2X1 U8064 ( .A(D3[4]), .B(in_valid), .Y(N5392) );
  AND2X1 U8065 ( .A(D3[3]), .B(in_valid), .Y(N5391) );
  AND2X1 U8066 ( .A(D3[2]), .B(in_valid), .Y(N5390) );
  AND2X1 U8067 ( .A(D3[1]), .B(in_valid), .Y(N5389) );
  AND2X1 U8068 ( .A(D3[0]), .B(in_valid), .Y(N5388) );
  AOI221XL U8069 ( .A0(y_out_sum11[9]), .A1(n364), .B0(y_out_sum11[8]), .B1(
        n365), .C0(n374), .Y(n373) );
  OAI22X1 U8070 ( .A0(n361), .A1(n4908), .B0(n359), .B1(n4856), .Y(n374) );
  AOI221XL U8071 ( .A0(y_out_sum8[9]), .A1(n421), .B0(y_out_sum8[8]), .B1(n422), .C0(n431), .Y(n430) );
  OAI22X1 U8072 ( .A0(n418), .A1(n4915), .B0(n416), .B1(n4864), .Y(n431) );
  NOR3BX1 U8073 ( .AN(n2525), .B(next[2]), .C(n4849), .Y(n2526) );
  INVX2 U8074 ( .A(shift[3]), .Y(n7531) );
  OAI2BB1X1 U8075 ( .A0N(N5767), .A1N(n4991), .B0(n6134), .Y(n3723) );
  INVX2 U8076 ( .A(matrix), .Y(n7192) );
  OAI2BB1X1 U8077 ( .A0N(N5685), .A1N(n4998), .B0(n6231), .Y(n3833) );
  OAI2BB1X1 U8078 ( .A0N(N5726), .A1N(n4989), .B0(n6182), .Y(n3778) );
  OAI2BB1X1 U8079 ( .A0N(N5808), .A1N(n4990), .B0(n6086), .Y(n3668) );
  NAND3X1 U8080 ( .A(next[1]), .B(next[0]), .C(n2526), .Y(n800) );
  OAI2BB1X1 U8081 ( .A0N(N5422), .A1N(n5005), .B0(n5945), .Y(n3974) );
  NOR2X1 U8082 ( .A(in_valid2), .B(in_valid), .Y(n4030) );
  NOR2X1 U8083 ( .A(n7270), .B(next[0]), .Y(n2524) );
  INVX2 U8084 ( .A(next[1]), .Y(n7270) );
  BUFX2 U8085 ( .A(n203), .Y(n5361) );
  NAND4X1 U8086 ( .A(shift[3]), .B(n7258), .C(n925), .D(n7530), .Y(n203) );
  BUFX2 U8087 ( .A(n205), .Y(n5362) );
  NAND4BX1 U8088 ( .AN(shift[5]), .B(n923), .C(shift[4]), .D(n7258), .Y(n205)
         );
  AOI22X1 U8089 ( .A0(N7874), .A1(n388), .B0(n389), .B1(n7561), .Y(n351) );
  OAI22X1 U8090 ( .A0(n390), .A1(n7560), .B0(N7873), .B1(n391), .Y(n389) );
  OAI22X1 U8091 ( .A0(n398), .A1(n7560), .B0(N7873), .B1(n399), .Y(n388) );
  AOI221XL U8092 ( .A0(y_out_sum11[17]), .A1(n364), .B0(y_out_sum11[16]), .B1(
        n365), .C0(n392), .Y(n391) );
  AOI221XL U8093 ( .A0(y_out_sum11[26]), .A1(n6923), .B0(y_out_sum11[27]), 
        .B1(n6932), .C0(n6919), .Y(n399) );
  OAI22X1 U8094 ( .A0(n6936), .A1(n6918), .B0(n6934), .B1(n6917), .Y(n6919) );
  AOI22X1 U8095 ( .A0(N7766), .A1(n445), .B0(n446), .B1(n7589), .Y(n408) );
  OAI22X1 U8096 ( .A0(n447), .A1(n7588), .B0(N7765), .B1(n448), .Y(n446) );
  OAI22X1 U8097 ( .A0(n455), .A1(n7588), .B0(N7765), .B1(n456), .Y(n445) );
  AOI221XL U8098 ( .A0(y_out_sum8[17]), .A1(n421), .B0(y_out_sum8[16]), .B1(
        n422), .C0(n449), .Y(n448) );
  AOI221XL U8099 ( .A0(y_out_sum8[26]), .A1(n6899), .B0(y_out_sum8[27]), .B1(
        n6908), .C0(n6895), .Y(n456) );
  OAI22X1 U8100 ( .A0(n6912), .A1(n6894), .B0(n6910), .B1(n6893), .Y(n6895) );
  XOR2X1 U8101 ( .A(reg_length14[5]), .B(n5017), .Y(n5016) );
  OR2X1 U8102 ( .A(reg_length14[4]), .B(n7111), .Y(n5017) );
  AOI221XL U8103 ( .A0(y_out_sum11[22]), .A1(n6923), .B0(y_out_sum11[23]), 
        .B1(n6932), .C0(n6922), .Y(n390) );
  OAI22X1 U8104 ( .A0(n6936), .A1(n6921), .B0(n6934), .B1(n6920), .Y(n6922) );
  AOI221XL U8105 ( .A0(y_out_sum8[22]), .A1(n6899), .B0(y_out_sum8[23]), .B1(
        n6908), .C0(n6898), .Y(n447) );
  OAI22X1 U8106 ( .A0(n6912), .A1(n6897), .B0(n6910), .B1(n6896), .Y(n6898) );
  NAND4X1 U8107 ( .A(shift[5]), .B(n7258), .C(n923), .D(n7532), .Y(n193) );
  AOI221XL U8108 ( .A0(y_out_sum11[30]), .A1(n6923), .B0(y_out_sum11[31]), 
        .B1(n6932), .C0(n6916), .Y(n398) );
  OAI22X1 U8109 ( .A0(n6936), .A1(n6915), .B0(n6934), .B1(n6914), .Y(n6916) );
  AOI221XL U8110 ( .A0(y_out_sum8[30]), .A1(n6899), .B0(y_out_sum8[31]), .B1(
        n6908), .C0(n6892), .Y(n455) );
  OAI22X1 U8111 ( .A0(n6912), .A1(n6891), .B0(n6910), .B1(n6890), .Y(n6892) );
  NAND3X1 U8112 ( .A(next[0]), .B(n7291), .C(next[1]), .Y(n745) );
  NOR2X1 U8113 ( .A(reg_length8[0]), .B(N7764), .Y(n421) );
  NOR2X1 U8114 ( .A(reg_length11[0]), .B(N7872), .Y(n364) );
  NOR2X1 U8115 ( .A(n5898), .B(next[1]), .Y(n2520) );
  NAND2X1 U8116 ( .A(N7944), .B(reg_length13[0]), .Y(n612) );
  OAI221X1 U8117 ( .A0(n592), .A1(n7538), .B0(n594), .B1(n7539), .C0(n596), 
        .Y(n582) );
  AOI222XL U8118 ( .A0(reg_length14[1]), .A1(n597), .B0(n598), .B1(n599), .C0(
        n600), .C1(n601), .Y(n596) );
  OAI222X1 U8119 ( .A0(n658), .A1(n7553), .B0(N7911), .B1(n660), .C0(n661), 
        .C1(n5024), .Y(n599) );
  OAI222X1 U8120 ( .A0(n602), .A1(n7545), .B0(N7947), .B1(n604), .C0(n605), 
        .C1(n5022), .Y(n601) );
  AOI221XL U8121 ( .A0(y_out_sum13[5]), .A1(n615), .B0(y_out_sum13[4]), .B1(
        n616), .C0(n636), .Y(n6829) );
  OAI22X1 U8122 ( .A0(n612), .A1(n4930), .B0(n610), .B1(n4874), .Y(n636) );
  AOI32X1 U8123 ( .A0(n7544), .A1(n5022), .A2(n621), .B0(N7946), .B1(n622), 
        .Y(n604) );
  OAI22X1 U8124 ( .A0(n623), .A1(n7543), .B0(N7945), .B1(n624), .Y(n622) );
  OAI22X1 U8125 ( .A0(N7945), .A1(n6830), .B0(n7543), .B1(n6829), .Y(n621) );
  AOI221XL U8126 ( .A0(y_out_sum13[13]), .A1(n615), .B0(y_out_sum13[12]), .B1(
        n616), .C0(n628), .Y(n623) );
  AOI221XL U8127 ( .A0(y_out_sum13[1]), .A1(n615), .B0(y_out_sum13[0]), .B1(
        n616), .C0(n6828), .Y(n6830) );
  OAI22X1 U8128 ( .A0(n610), .A1(n4880), .B0(n612), .B1(n4927), .Y(n6828) );
  AOI221XL U8129 ( .A0(y_out_sum13[9]), .A1(n615), .B0(y_out_sum13[8]), .B1(
        n616), .C0(n625), .Y(n624) );
  OAI22X1 U8130 ( .A0(n612), .A1(n4939), .B0(n610), .B1(n4886), .Y(n625) );
  INVX2 U8131 ( .A(shift[2]), .Y(n7530) );
  NAND2X1 U8132 ( .A(N7800), .B(reg_length9[0]), .Y(n534) );
  AOI221XL U8133 ( .A0(y_out_sum9[5]), .A1(n537), .B0(y_out_sum9[4]), .B1(n538), .C0(n558), .Y(n6853) );
  OAI22X1 U8134 ( .A0(n534), .A1(n4923), .B0(n532), .B1(n4871), .Y(n558) );
  AOI32X1 U8135 ( .A0(n7580), .A1(n5028), .A2(n543), .B0(N7802), .B1(n544), 
        .Y(n526) );
  OAI22X1 U8136 ( .A0(n545), .A1(n7579), .B0(N7801), .B1(n546), .Y(n544) );
  OAI22X1 U8137 ( .A0(N7801), .A1(n6854), .B0(n7579), .B1(n6853), .Y(n543) );
  AOI221XL U8138 ( .A0(y_out_sum9[13]), .A1(n537), .B0(y_out_sum9[12]), .B1(
        n538), .C0(n550), .Y(n545) );
  NAND2X1 U8139 ( .A(N7728), .B(reg_length7[0]), .Y(n478) );
  AOI221XL U8140 ( .A0(y_out_sum7[5]), .A1(n481), .B0(y_out_sum7[4]), .B1(n482), .C0(n502), .Y(n6877) );
  OAI22X1 U8141 ( .A0(n478), .A1(n4917), .B0(n476), .B1(n4867), .Y(n502) );
  AOI32X1 U8142 ( .A0(n7598), .A1(n5026), .A2(n487), .B0(N7730), .B1(n488), 
        .Y(n470) );
  OAI22X1 U8143 ( .A0(n489), .A1(n7597), .B0(N7729), .B1(n490), .Y(n488) );
  OAI22X1 U8144 ( .A0(N7729), .A1(n6878), .B0(n7597), .B1(n6877), .Y(n487) );
  AOI221XL U8145 ( .A0(y_out_sum7[13]), .A1(n481), .B0(y_out_sum7[12]), .B1(
        n482), .C0(n494), .Y(n489) );
  XOR2X1 U8146 ( .A(reg_length8[5]), .B(n5019), .Y(n5018) );
  OR2X1 U8147 ( .A(reg_length8[4]), .B(n7086), .Y(n5019) );
  INVX2 U8148 ( .A(shift[4]), .Y(n7532) );
  XOR2X1 U8149 ( .A(reg_length11[5]), .B(n5021), .Y(n5020) );
  OR2X1 U8150 ( .A(reg_length11[4]), .B(n7099), .Y(n5021) );
  AOI221XL U8151 ( .A0(y_out_sum9[1]), .A1(n537), .B0(y_out_sum9[0]), .B1(n538), .C0(n6852), .Y(n6854) );
  OAI22X1 U8152 ( .A0(n532), .A1(n4877), .B0(n534), .B1(n4922), .Y(n6852) );
  AOI221XL U8153 ( .A0(y_out_sum7[1]), .A1(n481), .B0(y_out_sum7[0]), .B1(n482), .C0(n6876), .Y(n6878) );
  OAI22X1 U8154 ( .A0(n476), .A1(n4869), .B0(n478), .B1(n4918), .Y(n6876) );
  AOI22X1 U8155 ( .A0(N7981), .A1(n292), .B0(n293), .B1(n7534), .Y(n290) );
  OAI221X1 U8156 ( .A0(n6960), .A1(n6954), .B0(n6958), .B1(n6953), .C0(n6952), 
        .Y(n292) );
  OAI221X1 U8157 ( .A0(n6961), .A1(n6960), .B0(n6959), .B1(n6958), .C0(n6957), 
        .Y(n293) );
  AOI2BB2X1 U8158 ( .B0(y_out_sum14[39]), .B1(n6956), .A0N(n297), .A1N(n6951), 
        .Y(n6952) );
  AOI2BB2X1 U8159 ( .B0(y_out_sum14[35]), .B1(n6956), .A0N(n297), .A1N(n6955), 
        .Y(n6957) );
  OAI2BB1X1 U8160 ( .A0N(N6418), .A1N(n4992), .B0(n6438), .Y(n3284) );
  OR2X1 U8161 ( .A(n6437), .B(n6441), .Y(n6438) );
  INVX2 U8162 ( .A(y_out_sum13[1]), .Y(n6437) );
  NOR2X1 U8163 ( .A(next[0]), .B(next[1]), .Y(n2493) );
  AOI221XL U8164 ( .A0(y_out_sum10[5]), .A1(n224), .B0(y_out_sum10[4]), .B1(
        n225), .C0(n239), .Y(n6982) );
  OAI22X1 U8165 ( .A0(n227), .A1(n4921), .B0(n229), .B1(n4868), .Y(n239) );
  AOI21X1 U8166 ( .A0(N7840), .A1(n212), .B0(n213), .Y(n194) );
  OAI22X1 U8167 ( .A0(N7837), .A1(n260), .B0(n261), .B1(n7569), .Y(n212) );
  OAI22X1 U8168 ( .A0(n214), .A1(n7572), .B0(N7839), .B1(n216), .Y(n213) );
  AOI221XL U8169 ( .A0(y_out_sum10[38]), .A1(n6980), .B0(y_out_sum10[39]), 
        .B1(n6979), .C0(n6967), .Y(n261) );
  AOI32X1 U8170 ( .A0(n7570), .A1(n7571), .A2(n219), .B0(N7838), .B1(n220), 
        .Y(n216) );
  OAI22X1 U8171 ( .A0(n221), .A1(n7569), .B0(N7837), .B1(n223), .Y(n220) );
  OAI22X1 U8172 ( .A0(N7837), .A1(n6983), .B0(n7569), .B1(n6982), .Y(n219) );
  AOI221XL U8173 ( .A0(y_out_sum10[13]), .A1(n224), .B0(y_out_sum10[12]), .B1(
        n225), .C0(n231), .Y(n221) );
  BUFX2 U8174 ( .A(reg_length10[0]), .Y(n5364) );
  AOI221XL U8175 ( .A0(y_out_sum12[5]), .A1(n671), .B0(y_out_sum12[4]), .B1(
        n672), .C0(n692), .Y(n6805) );
  OAI22X1 U8176 ( .A0(n668), .A1(n4937), .B0(n666), .B1(n4883), .Y(n692) );
  BUFX2 U8177 ( .A(reg_length12[0]), .Y(n5365) );
  AOI32X1 U8178 ( .A0(n7552), .A1(n5024), .A2(n677), .B0(N7910), .B1(n678), 
        .Y(n660) );
  OAI22X1 U8179 ( .A0(n679), .A1(n7551), .B0(N7909), .B1(n680), .Y(n678) );
  OAI22X1 U8180 ( .A0(N7909), .A1(n6806), .B0(n7551), .B1(n6805), .Y(n677) );
  AOI221XL U8181 ( .A0(y_out_sum12[13]), .A1(n671), .B0(y_out_sum12[12]), .B1(
        n672), .C0(n684), .Y(n679) );
  AOI221XL U8182 ( .A0(n224), .A1(y_out_sum10[1]), .B0(n225), .B1(
        y_out_sum10[0]), .C0(n6981), .Y(n6983) );
  OAI22X1 U8183 ( .A0(n229), .A1(n4870), .B0(n227), .B1(n4920), .Y(n6981) );
  AOI221XL U8184 ( .A0(y_out_sum9[9]), .A1(n537), .B0(y_out_sum9[8]), .B1(n538), .C0(n547), .Y(n546) );
  OAI22X1 U8185 ( .A0(n534), .A1(n4932), .B0(n532), .B1(n4881), .Y(n547) );
  AOI221XL U8186 ( .A0(y_out_sum7[9]), .A1(n481), .B0(y_out_sum7[8]), .B1(n482), .C0(n491), .Y(n490) );
  OAI22X1 U8187 ( .A0(n478), .A1(n4926), .B0(n476), .B1(n4875), .Y(n491) );
  AOI221XL U8188 ( .A0(y_out_sum12[1]), .A1(n671), .B0(y_out_sum12[0]), .B1(
        n672), .C0(n6804), .Y(n6806) );
  OAI22X1 U8189 ( .A0(n666), .A1(n4887), .B0(n668), .B1(n4933), .Y(n6804) );
  AOI22X1 U8190 ( .A0(N7946), .A1(n639), .B0(n640), .B1(n7544), .Y(n602) );
  OAI22X1 U8191 ( .A0(n641), .A1(n7543), .B0(N7945), .B1(n642), .Y(n640) );
  OAI22X1 U8192 ( .A0(n649), .A1(n7543), .B0(N7945), .B1(n650), .Y(n639) );
  AOI221XL U8193 ( .A0(y_out_sum13[17]), .A1(n615), .B0(y_out_sum13[16]), .B1(
        n616), .C0(n643), .Y(n642) );
  AOI221XL U8194 ( .A0(y_out_sum13[26]), .A1(n6827), .B0(y_out_sum13[27]), 
        .B1(n6836), .C0(n6823), .Y(n650) );
  OAI22X1 U8195 ( .A0(n6840), .A1(n6822), .B0(n6838), .B1(n6821), .Y(n6823) );
  AOI222XL U8196 ( .A0(temp_w_mat_idx[3]), .A1(n2590), .B0(temp_w_mat_idx[1]), 
        .B1(n2579), .C0(temp_w_mat_idx[2]), .C1(n2591), .Y(n2589) );
  AOI222XL U8197 ( .A0(temp_w_mat_idx[2]), .A1(n2590), .B0(temp_w_mat_idx[0]), 
        .B1(n2579), .C0(temp_w_mat_idx[1]), .C1(n2591), .Y(n2600) );
  AOI221XL U8198 ( .A0(y_out_sum13[22]), .A1(n6827), .B0(y_out_sum13[23]), 
        .B1(n6836), .C0(n6826), .Y(n641) );
  OAI22X1 U8199 ( .A0(n6840), .A1(n6825), .B0(n6838), .B1(n6824), .Y(n6826) );
  AOI221XL U8200 ( .A0(y_out_sum13[30]), .A1(n6827), .B0(y_out_sum13[31]), 
        .B1(n6836), .C0(n6820), .Y(n649) );
  OAI22X1 U8201 ( .A0(n6840), .A1(n6819), .B0(n6838), .B1(n6818), .Y(n6820) );
  AOI221XL U8202 ( .A0(y_out_sum10[9]), .A1(n224), .B0(y_out_sum10[8]), .B1(
        n225), .C0(n226), .Y(n223) );
  OAI22X1 U8203 ( .A0(n227), .A1(n4928), .B0(n229), .B1(n4876), .Y(n226) );
  NOR2X1 U8204 ( .A(reg_length13[0]), .B(N7944), .Y(n615) );
  AOI221XL U8205 ( .A0(y_out_sum12[9]), .A1(n671), .B0(y_out_sum12[8]), .B1(
        n672), .C0(n681), .Y(n680) );
  OAI22X1 U8206 ( .A0(n668), .A1(n4942), .B0(n666), .B1(n4890), .Y(n681) );
  AOI22X1 U8207 ( .A0(N7730), .A1(n505), .B0(n506), .B1(n7598), .Y(n468) );
  OAI22X1 U8208 ( .A0(n507), .A1(n7597), .B0(N7729), .B1(n508), .Y(n506) );
  OAI22X1 U8209 ( .A0(n515), .A1(n7597), .B0(N7729), .B1(n516), .Y(n505) );
  AOI221XL U8210 ( .A0(y_out_sum7[17]), .A1(n481), .B0(y_out_sum7[16]), .B1(
        n482), .C0(n509), .Y(n508) );
  AOI221XL U8211 ( .A0(y_out_sum7[26]), .A1(n6875), .B0(y_out_sum7[27]), .B1(
        n6884), .C0(n6871), .Y(n516) );
  OAI22X1 U8212 ( .A0(n6888), .A1(n6870), .B0(n6886), .B1(n6869), .Y(n6871) );
  AOI22X1 U8213 ( .A0(n356), .A1(n7560), .B0(N7873), .B1(n358), .Y(n354) );
  OAI221X1 U8214 ( .A0(n6936), .A1(n6930), .B0(n6934), .B1(n6929), .C0(n6928), 
        .Y(n356) );
  OAI221X1 U8215 ( .A0(n6937), .A1(n6936), .B0(n6935), .B1(n6934), .C0(n6933), 
        .Y(n358) );
  AOI2BB2X1 U8216 ( .B0(y_out_sum11[35]), .B1(n6932), .A0N(n361), .A1N(n6927), 
        .Y(n6928) );
  AOI2BB2X1 U8217 ( .B0(y_out_sum11[39]), .B1(n6932), .A0N(n361), .A1N(n6931), 
        .Y(n6933) );
  AOI221XL U8218 ( .A0(y_out_sum7[22]), .A1(n6875), .B0(y_out_sum7[23]), .B1(
        n6884), .C0(n6874), .Y(n507) );
  OAI22X1 U8219 ( .A0(n6888), .A1(n6873), .B0(n6886), .B1(n6872), .Y(n6874) );
  AOI22X1 U8220 ( .A0(n413), .A1(n7588), .B0(N7765), .B1(n415), .Y(n411) );
  OAI221X1 U8221 ( .A0(n6912), .A1(n6906), .B0(n6910), .B1(n6905), .C0(n6904), 
        .Y(n413) );
  OAI221X1 U8222 ( .A0(n6913), .A1(n6912), .B0(n6911), .B1(n6910), .C0(n6909), 
        .Y(n415) );
  AOI2BB2X1 U8223 ( .B0(y_out_sum8[35]), .B1(n6908), .A0N(n418), .A1N(n6903), 
        .Y(n6904) );
  AOI2BB2X1 U8224 ( .B0(y_out_sum8[39]), .B1(n6908), .A0N(n418), .A1N(n6907), 
        .Y(n6909) );
  AOI22X1 U8225 ( .A0(N7802), .A1(n561), .B0(n562), .B1(n7580), .Y(n524) );
  OAI22X1 U8226 ( .A0(n563), .A1(n7579), .B0(N7801), .B1(n564), .Y(n562) );
  OAI22X1 U8227 ( .A0(n571), .A1(n7579), .B0(N7801), .B1(n572), .Y(n561) );
  AOI221XL U8228 ( .A0(y_out_sum9[17]), .A1(n537), .B0(y_out_sum9[16]), .B1(
        n538), .C0(n565), .Y(n564) );
  AOI221XL U8229 ( .A0(y_out_sum9[26]), .A1(n6851), .B0(y_out_sum9[27]), .B1(
        n6860), .C0(n6847), .Y(n572) );
  OAI22X1 U8230 ( .A0(n6864), .A1(n6846), .B0(n6862), .B1(n6845), .Y(n6847) );
  OAI2BB1X1 U8231 ( .A0N(N5725), .A1N(n4989), .B0(n6184), .Y(n3779) );
  OR2X1 U8232 ( .A(n6186), .B(n6183), .Y(n6184) );
  INVX2 U8233 ( .A(y_out_sum4[1]), .Y(n6183) );
  OAI2BB1X1 U8234 ( .A0N(N5766), .A1N(n4991), .B0(n6136), .Y(n3724) );
  OR2X1 U8235 ( .A(n6138), .B(n6135), .Y(n6136) );
  INVX2 U8236 ( .A(y_out_sum5[1]), .Y(n6135) );
  OAI2BB1X1 U8237 ( .A0N(N5807), .A1N(n4990), .B0(n6088), .Y(n3669) );
  OR2X1 U8238 ( .A(n6090), .B(n6087), .Y(n6088) );
  INVX2 U8239 ( .A(y_out_sum6[1]), .Y(n6087) );
  OAI2BB1X1 U8240 ( .A0N(N6172), .A1N(n4994), .B0(n6768), .Y(n3614) );
  OR2X1 U8241 ( .A(n6767), .B(n6771), .Y(n6768) );
  INVX2 U8242 ( .A(y_out_sum7[1]), .Y(n6767) );
  OAI2BB1X1 U8243 ( .A0N(N6336), .A1N(n4999), .B0(n6546), .Y(n3394) );
  OR2X1 U8244 ( .A(n6545), .B(n6549), .Y(n6546) );
  INVX2 U8245 ( .A(y_out_sum11[1]), .Y(n6545) );
  OAI2BB1X1 U8246 ( .A0N(N6377), .A1N(n5000), .B0(n6492), .Y(n3339) );
  OR2X1 U8247 ( .A(n6491), .B(n6495), .Y(n6492) );
  INVX2 U8248 ( .A(y_out_sum12[1]), .Y(n6491) );
  OAI2BB1X1 U8249 ( .A0N(N6213), .A1N(n4995), .B0(n6713), .Y(n3559) );
  OR2X1 U8250 ( .A(n6712), .B(n6716), .Y(n6713) );
  INVX2 U8251 ( .A(y_out_sum8[1]), .Y(n6712) );
  OAI2BB1X1 U8252 ( .A0N(N6254), .A1N(n4996), .B0(n6658), .Y(n3504) );
  OR2X1 U8253 ( .A(n6657), .B(n6661), .Y(n6658) );
  INVX2 U8254 ( .A(y_out_sum9[1]), .Y(n6657) );
  OAI2BB1X1 U8255 ( .A0N(N6295), .A1N(n4997), .B0(n6602), .Y(n3449) );
  OR2X1 U8256 ( .A(n6601), .B(n6605), .Y(n6602) );
  INVX2 U8257 ( .A(y_out_sum10[1]), .Y(n6601) );
  OAI2BB1X1 U8258 ( .A0N(N6459), .A1N(n4993), .B0(n6384), .Y(n3229) );
  OR2X1 U8259 ( .A(n6383), .B(n6387), .Y(n6384) );
  INVX2 U8260 ( .A(y_out_sum14[1]), .Y(n6383) );
  OAI2BB1X1 U8261 ( .A0N(N5421), .A1N(n5005), .B0(n5947), .Y(n3975) );
  OR2X1 U8262 ( .A(n5949), .B(n5946), .Y(n5947) );
  INVX2 U8263 ( .A(y_out_sum0[1]), .Y(n5946) );
  AOI221XL U8264 ( .A0(y_out_sum7[30]), .A1(n6875), .B0(y_out_sum7[31]), .B1(
        n6884), .C0(n6868), .Y(n515) );
  OAI22X1 U8265 ( .A0(n6888), .A1(n6867), .B0(n6886), .B1(n6866), .Y(n6868) );
  AOI221XL U8266 ( .A0(y_out_sum9[22]), .A1(n6851), .B0(y_out_sum9[23]), .B1(
        n6860), .C0(n6850), .Y(n563) );
  OAI22X1 U8267 ( .A0(n6864), .A1(n6849), .B0(n6862), .B1(n6848), .Y(n6850) );
  OAI2BB1X1 U8268 ( .A0N(N5462), .A1N(n5003), .B0(n6334), .Y(n3935) );
  OR2X1 U8269 ( .A(n6336), .B(n6333), .Y(n6334) );
  INVX2 U8270 ( .A(y_out_sum1[1]), .Y(n6333) );
  OAI2BB1X1 U8271 ( .A0N(N5503), .A1N(n5002), .B0(n6284), .Y(n3889) );
  OR2X1 U8272 ( .A(n6286), .B(n6283), .Y(n6284) );
  INVX2 U8273 ( .A(y_out_sum2[1]), .Y(n6283) );
  OAI2BB1X1 U8274 ( .A0N(N5684), .A1N(n4998), .B0(n6233), .Y(n3834) );
  OR2X1 U8275 ( .A(n6235), .B(n6232), .Y(n6233) );
  INVX2 U8276 ( .A(y_out_sum3[1]), .Y(n6232) );
  AOI221XL U8277 ( .A0(y_out_sum9[30]), .A1(n6851), .B0(y_out_sum9[31]), .B1(
        n6860), .C0(n6844), .Y(n571) );
  OAI22X1 U8278 ( .A0(n6864), .A1(n6843), .B0(n6862), .B1(n6842), .Y(n6844) );
  NOR2X1 U8279 ( .A(reg_length9[0]), .B(N7800), .Y(n537) );
  NOR2X1 U8280 ( .A(reg_length7[0]), .B(N7728), .Y(n481) );
  AOI22X1 U8281 ( .A0(N7838), .A1(n242), .B0(n243), .B1(n7570), .Y(n214) );
  OAI22X1 U8282 ( .A0(n244), .A1(n7569), .B0(N7837), .B1(n245), .Y(n243) );
  OAI22X1 U8283 ( .A0(n252), .A1(n7569), .B0(N7837), .B1(n253), .Y(n242) );
  AOI221XL U8284 ( .A0(y_out_sum10[17]), .A1(n224), .B0(y_out_sum10[16]), .B1(
        n225), .C0(n246), .Y(n245) );
  AOI221XL U8285 ( .A0(y_out_sum10[26]), .A1(n6980), .B0(y_out_sum10[27]), 
        .B1(n6979), .C0(n6973), .Y(n253) );
  OAI22X1 U8286 ( .A0(n6977), .A1(n6972), .B0(n6975), .B1(n6971), .Y(n6973) );
  AOI22X1 U8287 ( .A0(N7910), .A1(n695), .B0(n696), .B1(n7552), .Y(n658) );
  OAI22X1 U8288 ( .A0(n697), .A1(n7551), .B0(N7909), .B1(n698), .Y(n696) );
  OAI22X1 U8289 ( .A0(n705), .A1(n7551), .B0(N7909), .B1(n706), .Y(n695) );
  AOI221XL U8290 ( .A0(y_out_sum12[17]), .A1(n671), .B0(y_out_sum12[16]), .B1(
        n672), .C0(n699), .Y(n698) );
  AOI221XL U8291 ( .A0(y_out_sum12[26]), .A1(n6803), .B0(y_out_sum12[27]), 
        .B1(n6812), .C0(n6799), .Y(n706) );
  OAI22X1 U8292 ( .A0(n6816), .A1(n6798), .B0(n6814), .B1(n6797), .Y(n6799) );
  INVX2 U8293 ( .A(count[1]), .Y(n7302) );
  AOI221XL U8294 ( .A0(y_out_sum10[22]), .A1(n6980), .B0(y_out_sum10[23]), 
        .B1(n6979), .C0(n6978), .Y(n244) );
  OAI22X1 U8295 ( .A0(n6977), .A1(n6976), .B0(n6975), .B1(n6974), .Y(n6978) );
  AOI221XL U8296 ( .A0(y_out_sum12[22]), .A1(n6803), .B0(y_out_sum12[23]), 
        .B1(n6812), .C0(n6802), .Y(n697) );
  OAI22X1 U8297 ( .A0(n6816), .A1(n6801), .B0(n6814), .B1(n6800), .Y(n6802) );
  AOI221XL U8298 ( .A0(y_out_sum10[30]), .A1(n6980), .B0(y_out_sum10[31]), 
        .B1(n6979), .C0(n6970), .Y(n252) );
  OAI22X1 U8299 ( .A0(n6977), .A1(n6969), .B0(n6975), .B1(n6968), .Y(n6970) );
  XOR2X1 U8300 ( .A(reg_length13[5]), .B(n5023), .Y(n5022) );
  OR2X1 U8301 ( .A(reg_length13[4]), .B(n7107), .Y(n5023) );
  AOI221XL U8302 ( .A0(y_out_sum12[30]), .A1(n6803), .B0(y_out_sum12[31]), 
        .B1(n6812), .C0(n6796), .Y(n705) );
  OAI22X1 U8303 ( .A0(n6816), .A1(n6795), .B0(n6814), .B1(n6794), .Y(n6796) );
  INVX2 U8304 ( .A(count[0]), .Y(n7303) );
  INVX2 U8305 ( .A(count[2]), .Y(n7304) );
  OAI2BB1X1 U8306 ( .A0N(reg_length0[3]), .A1N(n6005), .B0(n6033), .Y(N7432)
         );
  OR2X1 U8307 ( .A(reg_length0[1]), .B(reg_length0[0]), .Y(n6780) );
  OR2X1 U8308 ( .A(reg_length0[3]), .B(n6005), .Y(n6033) );
  OR2X1 U8309 ( .A(reg_length0[2]), .B(n6780), .Y(n6005) );
  INVX2 U8310 ( .A(count[3]), .Y(n7305) );
  XOR2X1 U8311 ( .A(reg_length12[5]), .B(n5025), .Y(n5024) );
  OR2X1 U8312 ( .A(reg_length12[4]), .B(n7103), .Y(n5025) );
  XOR2X1 U8313 ( .A(n5027), .B(n7081), .Y(n5026) );
  BUFX2 U8314 ( .A(N5058), .Y(n5379) );
  XOR2X1 U8315 ( .A(reg_length9[5]), .B(n5029), .Y(n5028) );
  OR2X1 U8316 ( .A(reg_length9[4]), .B(n7090), .Y(n5029) );
  OAI211X1 U8317 ( .A0(n170), .A1(n171), .B0(n580), .C0(n581), .Y(n6995) );
  AOI22X1 U8318 ( .A0(reg_length7[2]), .A1(n7255), .B0(reg_length7[1]), .B1(
        n7254), .Y(n170) );
  AOI221XL U8319 ( .A0(n714), .A1(reg_length7[4]), .B0(n715), .B1(
        reg_length7[5]), .C0(n7252), .Y(n581) );
  AOI211X1 U8320 ( .A0(n721), .A1(reg_length12[4]), .B0(n722), .C0(n7256), .Y(
        n580) );
  NAND2X1 U8321 ( .A(n754), .B(n755), .Y(n753) );
  AOI222XL U8322 ( .A0(reg_length4[1]), .A1(n7254), .B0(reg_length4[3]), .B1(
        n7257), .C0(reg_length4[2]), .C1(n7255), .Y(n754) );
  AOI222XL U8323 ( .A0(reg_length4[4]), .A1(n7244), .B0(reg_length4[0]), .B1(
        n7249), .C0(reg_length4[5]), .C1(n7260), .Y(n755) );
  OAI221X1 U8324 ( .A0(n897), .A1(n745), .B0(n7624), .B1(n761), .C0(n899), .Y(
        n837) );
  NOR4X1 U8325 ( .A(n913), .B(reg_length3[0]), .C(reg_length3[2]), .D(
        reg_length3[1]), .Y(n897) );
  INVX2 U8326 ( .A(n876), .Y(n7624) );
  AOI22X1 U8327 ( .A0(n7286), .A1(n900), .B0(n7277), .B1(n901), .Y(n899) );
  AOI22X1 U8328 ( .A0(n607), .A1(n7543), .B0(N7945), .B1(n609), .Y(n605) );
  OAI221X1 U8329 ( .A0(n6840), .A1(n6834), .B0(n6838), .B1(n6833), .C0(n6832), 
        .Y(n607) );
  OAI221X1 U8330 ( .A0(n6841), .A1(n6840), .B0(n6839), .B1(n6838), .C0(n6837), 
        .Y(n609) );
  AOI2BB2X1 U8331 ( .B0(y_out_sum13[35]), .B1(n6836), .A0N(n612), .A1N(n6831), 
        .Y(n6832) );
  AOI2BB2X1 U8332 ( .B0(y_out_sum13[39]), .B1(n6836), .A0N(n612), .A1N(n6835), 
        .Y(n6837) );
  BUFX2 U8333 ( .A(count[4]), .Y(n5380) );
  NAND2X1 U8334 ( .A(n756), .B(n757), .Y(n751) );
  AOI222XL U8335 ( .A0(reg_length6[1]), .A1(n7254), .B0(reg_length6[3]), .B1(
        n7257), .C0(reg_length6[2]), .C1(n7255), .Y(n756) );
  AOI222XL U8336 ( .A0(reg_length6[4]), .A1(n7244), .B0(reg_length6[0]), .B1(
        n7249), .C0(reg_length6[5]), .C1(n7260), .Y(n757) );
  AOI22X1 U8337 ( .A0(n529), .A1(n7579), .B0(N7801), .B1(n531), .Y(n527) );
  OAI221X1 U8338 ( .A0(n6864), .A1(n6858), .B0(n6862), .B1(n6857), .C0(n6856), 
        .Y(n529) );
  OAI221X1 U8339 ( .A0(n6865), .A1(n6864), .B0(n6863), .B1(n6862), .C0(n6861), 
        .Y(n531) );
  AOI2BB2X1 U8340 ( .B0(y_out_sum9[35]), .B1(n6860), .A0N(n534), .A1N(n6855), 
        .Y(n6856) );
  AOI222XL U8341 ( .A0(reg_length11[3]), .A1(n7257), .B0(reg_length11[5]), 
        .B1(n7260), .C0(reg_length11[4]), .C1(n7244), .Y(n207) );
  AOI221XL U8342 ( .A0(y_out_sum10[34]), .A1(n6980), .B0(y_out_sum10[35]), 
        .B1(n6979), .C0(n6964), .Y(n260) );
  OAI22X1 U8343 ( .A0(n6977), .A1(n6963), .B0(n6975), .B1(n6962), .Y(n6964) );
  OAI221X1 U8344 ( .A0(n6889), .A1(n6888), .B0(n6887), .B1(n6886), .C0(n6885), 
        .Y(n475) );
  AOI2BB2X1 U8345 ( .B0(y_out_sum7[39]), .B1(n6884), .A0N(n478), .A1N(n6883), 
        .Y(n6885) );
  NAND2X1 U8346 ( .A(n758), .B(n759), .Y(n749) );
  AOI222XL U8347 ( .A0(reg_length5[1]), .A1(n7254), .B0(reg_length5[3]), .B1(
        n7257), .C0(reg_length5[2]), .C1(n7255), .Y(n758) );
  AOI222XL U8348 ( .A0(reg_length5[4]), .A1(n7244), .B0(reg_length5[0]), .B1(
        n7249), .C0(reg_length5[5]), .C1(n7260), .Y(n759) );
  OAI2BB1X1 U8349 ( .A0N(reg_length0[1]), .A1N(reg_length0[0]), .B0(n6780), 
        .Y(N7430) );
  AOI22X1 U8350 ( .A0(n663), .A1(n7551), .B0(N7909), .B1(n665), .Y(n661) );
  OAI221X1 U8351 ( .A0(n6816), .A1(n6810), .B0(n6814), .B1(n6809), .C0(n6808), 
        .Y(n663) );
  OAI221X1 U8352 ( .A0(n6817), .A1(n6816), .B0(n6815), .B1(n6814), .C0(n6813), 
        .Y(n665) );
  AOI2BB2X1 U8353 ( .B0(y_out_sum12[35]), .B1(n6812), .A0N(n668), .A1N(n6807), 
        .Y(n6808) );
  AOI2BB2X1 U8354 ( .B0(y_out_sum12[39]), .B1(n6812), .A0N(n668), .A1N(n6811), 
        .Y(n6813) );
  OAI221X1 U8355 ( .A0(n6888), .A1(n6882), .B0(n6886), .B1(n6881), .C0(n6880), 
        .Y(n473) );
  AOI2BB2X1 U8356 ( .B0(y_out_sum7[35]), .B1(n6884), .A0N(n478), .A1N(n6879), 
        .Y(n6880) );
  OAI221X1 U8357 ( .A0(n7606), .A1(n1746), .B0(n5355), .B1(n7388), .C0(n1756), 
        .Y(n3619) );
  INVX2 U8358 ( .A(reg_length6[3]), .Y(n7606) );
  NAND2X1 U8359 ( .A(N7691), .B(n7218), .Y(n1756) );
  OAI221X1 U8360 ( .A0(n7608), .A1(n1746), .B0(n5355), .B1(n7392), .C0(n1749), 
        .Y(n3617) );
  INVX2 U8361 ( .A(reg_length6[5]), .Y(n7608) );
  NAND2X1 U8362 ( .A(N7693), .B(n7218), .Y(n1749) );
  OAI221X1 U8363 ( .A0(n7607), .A1(n1746), .B0(n5355), .B1(n7393), .C0(n1753), 
        .Y(n3618) );
  INVX2 U8364 ( .A(reg_length6[4]), .Y(n7607) );
  NAND2X1 U8365 ( .A(N7692), .B(n7218), .Y(n1753) );
  OAI211X1 U8366 ( .A0(n760), .A1(n761), .B0(n762), .C0(n763), .Y(n732) );
  AOI22X1 U8367 ( .A0(reg_length2[1]), .A1(n764), .B0(reg_length2[0]), .B1(
        n765), .Y(n763) );
  AOI221XL U8368 ( .A0(reg_length2[5]), .A1(n7260), .B0(reg_length2[4]), .B1(
        n7244), .C0(n768), .Y(n760) );
  OAI2BB1X1 U8369 ( .A0N(n766), .A1N(n767), .B0(n7285), .Y(n762) );
  AOI222XL U8370 ( .A0(reg_length1[4]), .A1(n7244), .B0(reg_length1[0]), .B1(
        n7249), .C0(reg_length1[5]), .C1(n7260), .Y(n767) );
  AOI222XL U8371 ( .A0(reg_length1[1]), .A1(n7254), .B0(reg_length1[3]), .B1(
        n7257), .C0(reg_length1[2]), .C1(n7255), .Y(n766) );
  OAI2BB1X1 U8372 ( .A0N(N5461), .A1N(n5003), .B0(n6337), .Y(n3936) );
  OR2X1 U8373 ( .A(n6336), .B(n6335), .Y(n6337) );
  INVX2 U8374 ( .A(y_out_sum1[0]), .Y(n6335) );
  OAI2BB1X1 U8375 ( .A0N(N5502), .A1N(n5002), .B0(n6287), .Y(n3890) );
  OR2X1 U8376 ( .A(n6286), .B(n6285), .Y(n6287) );
  INVX2 U8377 ( .A(y_out_sum2[0]), .Y(n6285) );
  OAI2BB1X1 U8378 ( .A0N(N5683), .A1N(n4998), .B0(n6236), .Y(n3835) );
  OR2X1 U8379 ( .A(n6235), .B(n6234), .Y(n6236) );
  INVX2 U8380 ( .A(y_out_sum3[0]), .Y(n6234) );
  OAI2BB1X1 U8381 ( .A0N(N5724), .A1N(n4989), .B0(n6187), .Y(n3780) );
  OR2X1 U8382 ( .A(n6186), .B(n6185), .Y(n6187) );
  INVX2 U8383 ( .A(y_out_sum4[0]), .Y(n6185) );
  OAI2BB1X1 U8384 ( .A0N(N5765), .A1N(n4991), .B0(n6139), .Y(n3725) );
  OR2X1 U8385 ( .A(n6138), .B(n6137), .Y(n6139) );
  INVX2 U8386 ( .A(y_out_sum5[0]), .Y(n6137) );
  OAI2BB1X1 U8387 ( .A0N(N5806), .A1N(n4990), .B0(n6091), .Y(n3670) );
  OR2X1 U8388 ( .A(n6090), .B(n6089), .Y(n6091) );
  INVX2 U8389 ( .A(y_out_sum6[0]), .Y(n6089) );
  OAI2BB1X1 U8390 ( .A0N(N6171), .A1N(n4994), .B0(n6770), .Y(n3615) );
  OR2X1 U8391 ( .A(n6769), .B(n6771), .Y(n6770) );
  INVX2 U8392 ( .A(y_out_sum7[0]), .Y(n6769) );
  OAI2BB1X1 U8393 ( .A0N(N6335), .A1N(n4999), .B0(n6548), .Y(n3395) );
  OR2X1 U8394 ( .A(n6547), .B(n6549), .Y(n6548) );
  INVX2 U8395 ( .A(y_out_sum11[0]), .Y(n6547) );
  OAI2BB1X1 U8396 ( .A0N(N5420), .A1N(n5005), .B0(n5950), .Y(n3976) );
  OR2X1 U8397 ( .A(n5949), .B(n5948), .Y(n5950) );
  INVX2 U8398 ( .A(y_out_sum0[0]), .Y(n5948) );
  OAI2BB1X1 U8399 ( .A0N(N6212), .A1N(n4995), .B0(n6715), .Y(n3560) );
  OR2X1 U8400 ( .A(n6714), .B(n6716), .Y(n6715) );
  INVX2 U8401 ( .A(y_out_sum8[0]), .Y(n6714) );
  OAI2BB1X1 U8402 ( .A0N(N6253), .A1N(n4996), .B0(n6660), .Y(n3505) );
  OR2X1 U8403 ( .A(n6659), .B(n6661), .Y(n6660) );
  INVX2 U8404 ( .A(y_out_sum9[0]), .Y(n6659) );
  OAI2BB1X1 U8405 ( .A0N(N6294), .A1N(n4997), .B0(n6604), .Y(n3450) );
  OR2X1 U8406 ( .A(n6603), .B(n6605), .Y(n6604) );
  INVX2 U8407 ( .A(y_out_sum10[0]), .Y(n6603) );
  OAI2BB1X1 U8408 ( .A0N(N6417), .A1N(n4992), .B0(n6440), .Y(n3285) );
  OR2X1 U8409 ( .A(n6439), .B(n6441), .Y(n6440) );
  INVX2 U8410 ( .A(y_out_sum13[0]), .Y(n6439) );
  XOR2X1 U8411 ( .A(n6033), .B(reg_length0[4]), .Y(n6032) );
  OAI2BB1X1 U8412 ( .A0N(N6376), .A1N(n5000), .B0(n6494), .Y(n3340) );
  OR2X1 U8413 ( .A(n6493), .B(n6495), .Y(n6494) );
  INVX2 U8414 ( .A(y_out_sum12[0]), .Y(n6493) );
  OAI2BB1X1 U8415 ( .A0N(N6458), .A1N(n4993), .B0(n6386), .Y(n3230) );
  OR2X1 U8416 ( .A(n6385), .B(n6387), .Y(n6386) );
  INVX2 U8417 ( .A(y_out_sum14[0]), .Y(n6385) );
  OAI222X1 U8418 ( .A0(n7551), .A1(n1435), .B0(n7555), .B1(n1436), .C0(n4850), 
        .C1(n7367), .Y(n3290) );
  INVX2 U8419 ( .A(reg_length12[2]), .Y(n7555) );
  OAI222X1 U8420 ( .A0(n7550), .A1(n1435), .B0(n7554), .B1(n1436), .C0(n4850), 
        .C1(n7366), .Y(n3291) );
  INVX2 U8421 ( .A(reg_length12[1]), .Y(n7554) );
  INVX2 U8422 ( .A(N7908), .Y(n7550) );
  OAI221X1 U8423 ( .A0(n7632), .A1(n2156), .B0(n5351), .B1(n7430), .C0(n2166), 
        .Y(n3894) );
  INVX2 U8424 ( .A(reg_length1[3]), .Y(n7632) );
  NAND2X1 U8425 ( .A(N7478), .B(n7209), .Y(n2166) );
  OAI221X1 U8426 ( .A0(n7634), .A1(n2156), .B0(n5351), .B1(n7434), .C0(n2159), 
        .Y(n3892) );
  INVX2 U8427 ( .A(reg_length1[5]), .Y(n7634) );
  NAND2X1 U8428 ( .A(N7480), .B(n7209), .Y(n2159) );
  OAI221X1 U8429 ( .A0(n7633), .A1(n2156), .B0(n5351), .B1(n7435), .C0(n2163), 
        .Y(n3893) );
  INVX2 U8430 ( .A(reg_length1[4]), .Y(n7633) );
  NAND2X1 U8431 ( .A(N7479), .B(n7209), .Y(n2163) );
  OAI222X1 U8432 ( .A0(n5022), .A1(n1381), .B0(n7549), .B1(n1383), .C0(n4847), 
        .C1(n7344), .Y(n3232) );
  INVX2 U8433 ( .A(reg_length13[5]), .Y(n7549) );
  OAI222X1 U8434 ( .A0(n7545), .A1(n1381), .B0(n7548), .B1(n1383), .C0(n4847), 
        .C1(n7345), .Y(n3233) );
  INVX2 U8435 ( .A(reg_length13[4]), .Y(n7548) );
  OAI222X1 U8436 ( .A0(n7544), .A1(n1381), .B0(n7547), .B1(n1383), .C0(n4847), 
        .C1(n7340), .Y(n3234) );
  INVX2 U8437 ( .A(reg_length13[3]), .Y(n7547) );
  OAI222X1 U8438 ( .A0(reg_length13[0]), .A1(n1381), .B0(N7943), .B1(n1383), 
        .C0(n4847), .C1(n7341), .Y(n3237) );
  XOR2X1 U8439 ( .A(n6034), .B(reg_length0[5]), .Y(n6040) );
  OR2X1 U8440 ( .A(reg_length0[4]), .B(n6033), .Y(n6034) );
  OAI221X1 U8441 ( .A0(n7619), .A1(n1994), .B0(n5353), .B1(n7412), .C0(n2008), 
        .Y(n3786) );
  INVX2 U8442 ( .A(reg_length3[1]), .Y(n7619) );
  NAND2X1 U8443 ( .A(N7566), .B(n7214), .Y(n2008) );
  OAI221X1 U8444 ( .A0(n7620), .A1(n1994), .B0(n5353), .B1(n7413), .C0(n2005), 
        .Y(n3785) );
  INVX2 U8445 ( .A(reg_length3[2]), .Y(n7620) );
  NAND2X1 U8446 ( .A(N7567), .B(n7214), .Y(n2005) );
  OAI222X1 U8447 ( .A0(reg_length9[0]), .A1(n1587), .B0(N7799), .B1(n1589), 
        .C0(n4851), .C1(n7353), .Y(n3457) );
  INVX2 U8448 ( .A(length9[0]), .Y(n7353) );
  INVX2 U8449 ( .A(length1[0]), .Y(n7431) );
  INVX2 U8450 ( .A(length6[0]), .Y(n7389) );
  INVX2 U8451 ( .A(length3[0]), .Y(n7411) );
  INVX2 U8452 ( .A(length2[0]), .Y(n7422) );
  INVX2 U8453 ( .A(length4[0]), .Y(n7403) );
  OAI222X1 U8454 ( .A0(reg_length11[0]), .A1(n1486), .B0(N7871), .B1(n1488), 
        .C0(n5359), .C1(n7371), .Y(n3347) );
  INVX2 U8455 ( .A(length11[0]), .Y(n7371) );
  INVX2 U8456 ( .A(length12[0]), .Y(n7365) );
  INVX2 U8457 ( .A(length13[0]), .Y(n7341) );
  INVX2 U8458 ( .A(length10[0]), .Y(n7347) );
  OAI222X1 U8459 ( .A0(n7599), .A1(n1691), .B0(n7603), .B1(n1693), .C0(n5356), 
        .C1(n7384), .Y(n3563) );
  INVX2 U8460 ( .A(reg_length7[4]), .Y(n7603) );
  OAI222X1 U8461 ( .A0(n7598), .A1(n1691), .B0(n7602), .B1(n1693), .C0(n5356), 
        .C1(n7379), .Y(n3564) );
  INVX2 U8462 ( .A(reg_length7[3]), .Y(n7602) );
  OAI222X1 U8463 ( .A0(reg_length7[0]), .A1(n1691), .B0(N7727), .B1(n1693), 
        .C0(n5356), .C1(n7380), .Y(n3567) );
  OAI222X1 U8464 ( .A0(n5020), .A1(n1486), .B0(n7567), .B1(n1488), .C0(n5359), 
        .C1(n7374), .Y(n3342) );
  INVX2 U8465 ( .A(reg_length11[5]), .Y(n7567) );
  OAI222X1 U8466 ( .A0(n7562), .A1(n1486), .B0(n7566), .B1(n1488), .C0(n5359), 
        .C1(n7375), .Y(n3343) );
  INVX2 U8467 ( .A(reg_length11[4]), .Y(n7566) );
  OAI222X1 U8468 ( .A0(n7561), .A1(n1486), .B0(n7565), .B1(n1488), .C0(n5359), 
        .C1(n7370), .Y(n3344) );
  INVX2 U8469 ( .A(reg_length11[3]), .Y(n7565) );
  AOI222XL U8470 ( .A0(reg_length3[4]), .A1(n7244), .B0(reg_length3[0]), .B1(
        n7249), .C0(reg_length3[5]), .C1(n7260), .Y(n772) );
  INVX2 U8471 ( .A(length7[0]), .Y(n7380) );
  OAI2BB2X1 U8472 ( .B0(n4851), .B1(n7353), .A0N(n7223), .A1N(reg_length09[0]), 
        .Y(n3466) );
  OAI2BB2X1 U8473 ( .B0(n5359), .B1(n7371), .A0N(n7225), .A1N(reg_length011[0]), .Y(n3356) );
  OAI2BB2X1 U8474 ( .B0(n4850), .B1(n7365), .A0N(n7226), .A1N(reg_length012[0]), .Y(n3301) );
  OAI2BB2X1 U8475 ( .B0(n4847), .B1(n7341), .A0N(n7227), .A1N(reg_length013[0]), .Y(n3246) );
  OAI2BB2X1 U8476 ( .B0(n5360), .B1(n7335), .A0N(n7228), .A1N(reg_length014[0]), .Y(n3191) );
  INVX2 U8477 ( .A(length14[0]), .Y(n7335) );
  OAI2BB2X1 U8478 ( .B0(n5358), .B1(n7347), .A0N(n7224), .A1N(reg_length010[0]), .Y(n3411) );
  AOI222XL U8479 ( .A0(reg_length3[1]), .A1(n7254), .B0(reg_length3[3]), .B1(
        n7257), .C0(reg_length3[2]), .C1(n7255), .Y(n771) );
  INVX2 U8480 ( .A(length5[0]), .Y(n7395) );
  INVX2 U8481 ( .A(y_out_sum11[24]), .Y(n6917) );
  OAI2BB2X1 U8482 ( .B0(n5356), .B1(n7380), .A0N(n7221), .A1N(reg_length07[0]), 
        .Y(n3576) );
  OAI2BB2X1 U8483 ( .B0(n5357), .B1(n7359), .A0N(n7222), .A1N(reg_length08[0]), 
        .Y(n3521) );
  INVX2 U8484 ( .A(length8[0]), .Y(n7359) );
  OAI2BB2X1 U8485 ( .B0(n5355), .B1(n7389), .A0N(n7219), .A1N(reg_length06[0]), 
        .Y(n3631) );
  OAI221X1 U8486 ( .A0(n7616), .A1(n1913), .B0(n5354), .B1(n7402), .C0(n1923), 
        .Y(n3729) );
  INVX2 U8487 ( .A(reg_length4[3]), .Y(n7616) );
  NAND2X1 U8488 ( .A(N7609), .B(n7216), .Y(n1923) );
  OAI222X1 U8489 ( .A0(reg_length14[0]), .A1(n1327), .B0(n4952), .B1(n1328), 
        .C0(n5360), .C1(n7335), .Y(n3182) );
  NAND4X1 U8490 ( .A(n7614), .B(n7615), .C(N7606), .D(n905), .Y(n901) );
  NOR3X1 U8491 ( .A(reg_length4[3]), .B(reg_length4[5]), .C(reg_length4[4]), 
        .Y(n905) );
  OAI221X1 U8492 ( .A0(n7618), .A1(n1913), .B0(n5354), .B1(n7406), .C0(n1916), 
        .Y(n3727) );
  INVX2 U8493 ( .A(reg_length4[5]), .Y(n7618) );
  NAND2X1 U8494 ( .A(N7611), .B(n7216), .Y(n1916) );
  OAI221X1 U8495 ( .A0(n7617), .A1(n1913), .B0(n5354), .B1(n7407), .C0(n1920), 
        .Y(n3728) );
  INVX2 U8496 ( .A(reg_length4[4]), .Y(n7617) );
  NAND2X1 U8497 ( .A(N7610), .B(n7216), .Y(n1920) );
  INVX2 U8498 ( .A(y_out_sum11[20]), .Y(n6920) );
  OAI222X1 U8499 ( .A0(reg_length8[0]), .A1(n1642), .B0(n4902), .B1(n1643), 
        .C0(n5357), .C1(n7359), .Y(n3512) );
  OAI222X1 U8500 ( .A0(n5026), .A1(n1691), .B0(n5027), .B1(n1693), .C0(n5356), 
        .C1(n7383), .Y(n3562) );
  INVX2 U8501 ( .A(y_out_sum14[24]), .Y(n6941) );
  INVX2 U8502 ( .A(y_out_sum11[25]), .Y(n6918) );
  INVX2 U8503 ( .A(N5060), .Y(n5572) );
  INVX2 U8504 ( .A(n717), .Y(n7252) );
  AOI222XL U8505 ( .A0(reg_length13[2]), .A1(n718), .B0(reg_length14[5]), .B1(
        n719), .C0(reg_length13[0]), .C1(n720), .Y(n717) );
  OAI2BB2X1 U8506 ( .B0(n5355), .B1(n7393), .A0N(n7219), .A1N(reg_length06[4]), 
        .Y(n3627) );
  OAI2BB2X1 U8507 ( .B0(n5355), .B1(n7388), .A0N(n7219), .A1N(reg_length06[3]), 
        .Y(n3628) );
  OAI2BB2X1 U8508 ( .B0(n5355), .B1(n7392), .A0N(n7219), .A1N(reg_length06[5]), 
        .Y(n3626) );
  INVX2 U8509 ( .A(y_out_sum14[20]), .Y(n6944) );
  OAI22X1 U8510 ( .A0(n2500), .A1(n2501), .B0(n2502), .B1(n2503), .Y(n2499) );
  NAND4X1 U8511 ( .A(n7626), .B(n7627), .C(n7628), .D(n7629), .Y(n2500) );
  NAND4X1 U8512 ( .A(n7610), .B(n7611), .C(n7612), .D(n7613), .Y(n2502) );
  NAND4X1 U8513 ( .A(reg_length5[0]), .B(n7286), .C(n2417), .D(n7609), .Y(
        n2503) );
  OAI2BB2X1 U8514 ( .B0(n2366), .B1(n7296), .A0N(N8524), .A1N(n7204), .Y(n4003) );
  INVX2 U8515 ( .A(next[7]), .Y(n7296) );
  OAI2BB2X1 U8516 ( .B0(n2366), .B1(n7295), .A0N(N8523), .A1N(n7204), .Y(n4004) );
  INVX2 U8517 ( .A(next[6]), .Y(n7295) );
  OAI2BB2X1 U8518 ( .B0(n2366), .B1(n7294), .A0N(N8522), .A1N(n7204), .Y(n4005) );
  INVX2 U8519 ( .A(next[5]), .Y(n7294) );
  OAI2BB2X1 U8520 ( .B0(n2366), .B1(n7293), .A0N(N8521), .A1N(n7204), .Y(n4006) );
  INVX2 U8521 ( .A(next[4]), .Y(n7293) );
  NAND4X1 U8522 ( .A(reg_length2[0]), .B(n7261), .C(n2413), .D(n7625), .Y(
        n2501) );
  AOI221XL U8523 ( .A0(n2495), .A1(n2496), .B0(n2497), .B1(n2498), .C0(n2499), 
        .Y(n2469) );
  NOR4X1 U8524 ( .A(reg_length3[5]), .B(reg_length3[4]), .C(reg_length3[3]), 
        .D(reg_length3[2]), .Y(n2496) );
  NOR4X1 U8525 ( .A(reg_length1[5]), .B(reg_length1[4]), .C(reg_length1[3]), 
        .D(reg_length1[2]), .Y(n2498) );
  NOR4X1 U8526 ( .A(reg_length1[1]), .B(n2420), .C(n802), .D(N7475), .Y(n2497)
         );
  NAND2X1 U8527 ( .A(n2389), .B(n2390), .Y(n2388) );
  OAI32X1 U8528 ( .A0(n2273), .A1(count1[0]), .A2(n2272), .B0(n2391), .B1(
        n5350), .Y(n2390) );
  NOR4X1 U8529 ( .A(n2392), .B(n2393), .C(n2394), .D(n2395), .Y(n2391) );
  NAND2X1 U8530 ( .A(n2399), .B(n2400), .Y(n2393) );
  NOR4X1 U8531 ( .A(reg_length7[1]), .B(n2514), .C(n171), .D(N7727), .Y(n2512)
         );
  NOR4X1 U8532 ( .A(n2515), .B(reg_length07[3]), .C(reg_length07[5]), .D(
        reg_length07[4]), .Y(n2514) );
  NAND3X1 U8533 ( .A(n4944), .B(n4892), .C(reg_length07[0]), .Y(n2515) );
  OAI2BB2X1 U8534 ( .B0(n5898), .B1(n2366), .A0N(N8517), .A1N(n7204), .Y(n4009) );
  INVX2 U8535 ( .A(y_out_sum14[25]), .Y(n6942) );
  NAND4X1 U8536 ( .A(n7609), .B(n7610), .C(n4934), .D(n909), .Y(n900) );
  NOR3X1 U8537 ( .A(reg_length5[3]), .B(reg_length5[5]), .C(reg_length5[4]), 
        .Y(n909) );
  INVX2 U8538 ( .A(y_out_sum11[21]), .Y(n6921) );
  INVX2 U8539 ( .A(N5059), .Y(n5573) );
  INVX2 U8540 ( .A(y_out_sum11[28]), .Y(n6914) );
  OAI2BB2X1 U8541 ( .B0(n5351), .B1(n7431), .A0N(n7210), .A1N(n2816), .Y(n3986) );
  OAI2BB2X1 U8542 ( .B0(n7197), .B1(n7395), .A0N(n7196), .A1N(n2820), .Y(n3686) );
  OAI2BB2X1 U8543 ( .B0(n5353), .B1(n7411), .A0N(n7215), .A1N(n2818), .Y(n3796) );
  OAI2BB2X1 U8544 ( .B0(n7213), .B1(n7422), .A0N(n7212), .A1N(n2817), .Y(n3851) );
  OAI2BB2X1 U8545 ( .B0(n5354), .B1(n7403), .A0N(n7217), .A1N(n2819), .Y(n3741) );
  INVX2 U8546 ( .A(y_out_sum14[21]), .Y(n6945) );
  AOI222XL U8547 ( .A0(reg_length8[2]), .A1(n589), .B0(reg_length7[3]), .B1(
        n590), .C0(reg_length8[1]), .C1(n591), .Y(n588) );
  OAI221X1 U8548 ( .A0(reg_invalid2[0]), .A1(n1484), .B0(n1864), .B1(n2800), 
        .C0(n2811), .Y(n2775) );
  AOI221XL U8549 ( .A0(n2700), .A1(n7046), .B0(n2716), .B1(n2710), .C0(n2727), 
        .Y(n2811) );
  INVX2 U8550 ( .A(y_out_sum14[28]), .Y(n6938) );
  NAND2X1 U8551 ( .A(n7285), .B(n891), .Y(n875) );
  NAND4X1 U8552 ( .A(n7630), .B(n7631), .C(N7475), .D(n895), .Y(n891) );
  NOR3X1 U8553 ( .A(reg_length1[3]), .B(reg_length1[5]), .C(reg_length1[4]), 
        .Y(n895) );
  INVX2 U8554 ( .A(y_out_sum11[29]), .Y(n6915) );
  OAI33X1 U8555 ( .A0(n7507), .A1(count12[0]), .A2(n1456), .B0(n1348), .B1(
        count14[0]), .B2(n7269), .Y(n2395) );
  INVX2 U8556 ( .A(length9[1]), .Y(n7354) );
  NAND4X1 U8557 ( .A(n5015), .B(n4944), .C(reg_length07[0]), .D(n2419), .Y(
        n1713) );
  NOR4X1 U8558 ( .A(reg_length07[5]), .B(reg_length07[4]), .C(reg_length07[3]), 
        .D(n2823), .Y(n2419) );
  INVX2 U8559 ( .A(y_out_sum14[29]), .Y(n6939) );
  OAI221X1 U8560 ( .A0(n94), .A1(n96), .B0(current_state[1]), .B1(n7194), .C0(
        n98), .Y(next_state[0]) );
  INVX2 U8561 ( .A(n93), .Y(n7194) );
  AOI31X1 U8562 ( .A0(n99), .A1(n7300), .A2(n101), .B0(n102), .Y(n98) );
  NOR4X1 U8563 ( .A(current_state[0]), .B(count[14]), .C(n5377), .D(N5118), 
        .Y(n101) );
  AND4X2 U8564 ( .A(count_state_idle[2]), .B(count_state_idle[1]), .C(
        count_state_idle[3]), .D(n123), .Y(n94) );
  NOR4X1 U8565 ( .A(n2858), .B(count_state_idle[5]), .C(count_state_idle[4]), 
        .D(n7033), .Y(n123) );
  OAI2BB2X1 U8566 ( .B0(n7197), .B1(n7398), .A0N(n7196), .A1N(reg_length05[5]), 
        .Y(n3681) );
  OAI2BB2X1 U8567 ( .B0(n7197), .B1(n7399), .A0N(n7196), .A1N(reg_length05[4]), 
        .Y(n3682) );
  OAI2BB2X1 U8568 ( .B0(n7197), .B1(n7394), .A0N(n7196), .A1N(reg_length05[3]), 
        .Y(n3683) );
  OAI2BB2X1 U8569 ( .B0(n5351), .B1(n7435), .A0N(n7210), .A1N(reg_length01[4]), 
        .Y(n3985) );
  OAI2BB2X1 U8570 ( .B0(n5351), .B1(n7430), .A0N(n7210), .A1N(reg_length01[3]), 
        .Y(n3984) );
  OAI2BB2X1 U8571 ( .B0(n5351), .B1(n7434), .A0N(n7210), .A1N(reg_length01[5]), 
        .Y(n4010) );
  AOI221XL U8572 ( .A0(reg_length11[0]), .A1(n7272), .B0(n5365), .B1(n7281), 
        .C0(n270), .Y(n192) );
  OAI22X1 U8573 ( .A0(n171), .A1(N7727), .B0(n272), .B1(n4902), .Y(n270) );
  NAND4X1 U8574 ( .A(n7625), .B(n7626), .C(N7521), .D(n912), .Y(n876) );
  NOR3X1 U8575 ( .A(reg_length2[3]), .B(reg_length2[5]), .C(reg_length2[4]), 
        .Y(n912) );
  OAI22X1 U8576 ( .A0(n2477), .A1(n2478), .B0(n2479), .B1(n2480), .Y(n2476) );
  NAND4X1 U8577 ( .A(n7583), .B(n7584), .C(n7585), .D(n7586), .Y(n2479) );
  NAND4X1 U8578 ( .A(n7574), .B(n7575), .C(n7576), .D(n7577), .Y(n2477) );
  NAND4X1 U8579 ( .A(reg_length9[0]), .B(n199), .C(n2402), .D(n7582), .Y(n2480) );
  INVX2 U8580 ( .A(y_out_sum8[24]), .Y(n6893) );
  INVX2 U8581 ( .A(y_out_sum8[20]), .Y(n6896) );
  OAI2BB2X1 U8582 ( .B0(n4850), .B1(n7369), .A0N(n7226), .A1N(reg_length012[4]), .Y(n3297) );
  OAI2BB2X1 U8583 ( .B0(n4850), .B1(n7368), .A0N(n7226), .A1N(reg_length012[5]), .Y(n3296) );
  OAI2BB2X1 U8584 ( .B0(n4850), .B1(n7364), .A0N(n7226), .A1N(reg_length012[3]), .Y(n3298) );
  INVX2 U8585 ( .A(length7[1]), .Y(n7381) );
  INVX2 U8586 ( .A(length11[1]), .Y(n7372) );
  INVX2 U8587 ( .A(length12[1]), .Y(n7366) );
  INVX2 U8588 ( .A(length8[1]), .Y(n7360) );
  INVX2 U8589 ( .A(length14[1]), .Y(n7336) );
  OAI2BB2X1 U8590 ( .B0(n5353), .B1(n7415), .A0N(n7215), .A1N(reg_length03[4]), 
        .Y(n3792) );
  OAI2BB2X1 U8591 ( .B0(n5353), .B1(n7410), .A0N(n7215), .A1N(reg_length03[3]), 
        .Y(n3793) );
  OAI2BB2X1 U8592 ( .B0(n5353), .B1(n7414), .A0N(n7215), .A1N(reg_length03[5]), 
        .Y(n3791) );
  INVX2 U8593 ( .A(y_out_sum8[25]), .Y(n6894) );
  INVX2 U8594 ( .A(length10[1]), .Y(n7348) );
  INVX2 U8595 ( .A(n142), .Y(n7200) );
  AOI22X1 U8596 ( .A0(count_state_idle[3]), .A1(n7203), .B0(N4524), .B1(n5350), 
        .Y(n142) );
  INVX2 U8597 ( .A(n143), .Y(n7201) );
  AOI22X1 U8598 ( .A0(count_state_idle[2]), .A1(n7203), .B0(N4523), .B1(n5350), 
        .Y(n143) );
  INVX2 U8599 ( .A(n144), .Y(n7202) );
  AOI22X1 U8600 ( .A0(count_state_idle[1]), .A1(n7203), .B0(N4522), .B1(n5350), 
        .Y(n144) );
  INVX2 U8601 ( .A(reg_length4[2]), .Y(n7615) );
  OAI2BB2X1 U8602 ( .B0(n4847), .B1(n7345), .A0N(n7227), .A1N(reg_length013[4]), .Y(n3242) );
  OAI2BB2X1 U8603 ( .B0(n4847), .B1(n7344), .A0N(n7227), .A1N(reg_length013[5]), .Y(n3241) );
  OAI2BB2X1 U8604 ( .B0(n4847), .B1(n7340), .A0N(n7227), .A1N(reg_length013[3]), .Y(n3243) );
  INVX2 U8605 ( .A(n141), .Y(n7199) );
  AOI22X1 U8606 ( .A0(n7203), .A1(count_state_idle[4]), .B0(N4525), .B1(n5350), 
        .Y(n141) );
  INVX2 U8607 ( .A(n138), .Y(n7198) );
  AOI22X1 U8608 ( .A0(n7203), .A1(count_state_idle[5]), .B0(N4526), .B1(n5350), 
        .Y(n138) );
  INVX2 U8609 ( .A(y_out_sum8[21]), .Y(n6897) );
  NOR4X1 U8610 ( .A(reg_length3[1]), .B(n2415), .C(n745), .D(N7565), .Y(n2495)
         );
  AOI211X1 U8611 ( .A0(n7267), .A1(n2466), .B0(n2467), .C0(n2394), .Y(n2465)
         );
  OAI32X1 U8612 ( .A0(n2521), .A1(n4952), .A2(n2522), .B0(count14[0]), .B1(
        n1348), .Y(n2466) );
  OAI33X1 U8613 ( .A0(n7507), .A1(count12[0]), .A2(n178), .B0(n1403), .B1(
        count13[0]), .B2(n169), .Y(n2467) );
  NAND4X1 U8614 ( .A(n7538), .B(n7539), .C(n7540), .D(n7541), .Y(n2521) );
  NAND4X1 U8615 ( .A(n7290), .B(n4945), .C(reg_length013[0]), .D(n2403), .Y(
        n1402) );
  NOR4X1 U8616 ( .A(reg_length013[5]), .B(reg_length013[4]), .C(
        reg_length013[3]), .D(n2835), .Y(n2403) );
  INVX2 U8617 ( .A(y_out_sum8[28]), .Y(n6890) );
  INVX2 U8618 ( .A(reg_length4[1]), .Y(n7614) );
  OAI2BB1X1 U8619 ( .A0N(reg_length0[2]), .A1N(n6780), .B0(n6005), .Y(N7431)
         );
  NAND4X1 U8620 ( .A(n7604), .B(n7605), .C(N7688), .D(n888), .Y(n836) );
  NOR3X1 U8621 ( .A(reg_length6[3]), .B(reg_length6[5]), .C(reg_length6[4]), 
        .Y(n888) );
  OAI2BB2X1 U8622 ( .B0(n7213), .B1(n7425), .A0N(n7212), .A1N(reg_length02[5]), 
        .Y(n3846) );
  OAI2BB2X1 U8623 ( .B0(n7213), .B1(n7426), .A0N(n7212), .A1N(reg_length02[4]), 
        .Y(n3847) );
  OAI2BB2X1 U8624 ( .B0(n7213), .B1(n7421), .A0N(n7212), .A1N(reg_length02[3]), 
        .Y(n3848) );
  NOR4X1 U8625 ( .A(reg_length8[1]), .B(n2418), .C(n272), .D(n4902), .Y(n2487)
         );
  NOR4X1 U8626 ( .A(reg_length4[1]), .B(n2414), .C(n867), .D(N7606), .Y(n2489)
         );
  INVX2 U8627 ( .A(length13[1]), .Y(n7342) );
  INVX2 U8628 ( .A(y_out_sum8[29]), .Y(n6891) );
  INVX2 U8629 ( .A(reg_length5[2]), .Y(n7610) );
  NOR4X1 U8630 ( .A(reg_length13[1]), .B(n2516), .C(n169), .D(N7943), .Y(n2510) );
  NOR4X1 U8631 ( .A(n2517), .B(reg_length013[3]), .C(reg_length013[5]), .D(
        reg_length013[4]), .Y(n2516) );
  NAND3X1 U8632 ( .A(n4945), .B(n4893), .C(reg_length013[0]), .Y(n2517) );
  NOR4X1 U8633 ( .A(reg_length12[1]), .B(n2398), .C(n178), .D(N7907), .Y(n2474) );
  INVX2 U8634 ( .A(reg_length5[1]), .Y(n7609) );
  OAI2BB2X1 U8635 ( .B0(n5354), .B1(n7407), .A0N(n7217), .A1N(reg_length04[4]), 
        .Y(n3737) );
  OAI2BB2X1 U8636 ( .B0(n5354), .B1(n7402), .A0N(n7217), .A1N(reg_length04[3]), 
        .Y(n3738) );
  OAI2BB2X1 U8637 ( .B0(n5354), .B1(n7406), .A0N(n7217), .A1N(reg_length04[5]), 
        .Y(n3736) );
  NAND4X1 U8638 ( .A(n7264), .B(n4948), .C(reg_length06[0]), .D(n2416), .Y(
        n1773) );
  NOR4X1 U8639 ( .A(reg_length06[5]), .B(reg_length06[4]), .C(reg_length06[3]), 
        .D(n2821), .Y(n2416) );
  OAI2BB2X1 U8640 ( .B0(n5358), .B1(n7351), .A0N(n7224), .A1N(reg_length010[4]), .Y(n3407) );
  OAI2BB2X1 U8641 ( .B0(n5358), .B1(n7346), .A0N(n7224), .A1N(reg_length010[3]), .Y(n3408) );
  OAI2BB2X1 U8642 ( .B0(n5358), .B1(n7350), .A0N(n7224), .A1N(reg_length010[5]), .Y(n3406) );
  OAI2BB2X1 U8643 ( .B0(n5356), .B1(n7384), .A0N(n7221), .A1N(reg_length07[4]), 
        .Y(n3572) );
  OAI2BB2X1 U8644 ( .B0(n5357), .B1(n7363), .A0N(n7222), .A1N(reg_length08[4]), 
        .Y(n3517) );
  OAI2BB2X1 U8645 ( .B0(n5356), .B1(n7383), .A0N(n7221), .A1N(reg_length07[5]), 
        .Y(n3571) );
  OAI2BB2X1 U8646 ( .B0(n5356), .B1(n7379), .A0N(n7221), .A1N(reg_length07[3]), 
        .Y(n3573) );
  OAI2BB2X1 U8647 ( .B0(n5357), .B1(n7362), .A0N(n7222), .A1N(reg_length08[5]), 
        .Y(n3516) );
  OAI2BB2X1 U8648 ( .B0(n5357), .B1(n7358), .A0N(n7222), .A1N(reg_length08[3]), 
        .Y(n3518) );
  INVX2 U8649 ( .A(reg_length3[3]), .Y(n7621) );
  OAI2BB2X1 U8650 ( .B0(n5360), .B1(n7339), .A0N(n7228), .A1N(reg_length014[4]), .Y(n3187) );
  OAI2BB2X1 U8651 ( .B0(n5360), .B1(n7338), .A0N(n7228), .A1N(reg_length014[5]), .Y(n3186) );
  OAI2BB2X1 U8652 ( .B0(n5360), .B1(n7334), .A0N(n7228), .A1N(reg_length014[3]), .Y(n3188) );
  OAI2BB2X1 U8653 ( .B0(n5359), .B1(n7375), .A0N(n7225), .A1N(reg_length011[4]), .Y(n3352) );
  OAI2BB2X1 U8654 ( .B0(n4851), .B1(n7357), .A0N(n7223), .A1N(reg_length09[4]), 
        .Y(n3462) );
  OAI2BB2X1 U8655 ( .B0(n5359), .B1(n7374), .A0N(n7225), .A1N(reg_length011[5]), .Y(n3351) );
  OAI2BB2X1 U8656 ( .B0(n5359), .B1(n7370), .A0N(n7225), .A1N(reg_length011[3]), .Y(n3353) );
  OAI2BB2X1 U8657 ( .B0(n4851), .B1(n7352), .A0N(n7223), .A1N(reg_length09[3]), 
        .Y(n3463) );
  OAI2BB2X1 U8658 ( .B0(n4851), .B1(n7356), .A0N(n7223), .A1N(reg_length09[5]), 
        .Y(n3461) );
  INVX2 U8659 ( .A(reg_length3[5]), .Y(n7623) );
  INVX2 U8660 ( .A(N5061), .Y(n5570) );
  INVX2 U8661 ( .A(reg_length3[4]), .Y(n7622) );
  INVX2 U8662 ( .A(N5062), .Y(n5569) );
  INVX2 U8663 ( .A(length1[1]), .Y(n7432) );
  INVX2 U8664 ( .A(length3[1]), .Y(n7412) );
  INVX2 U8665 ( .A(length5[1]), .Y(n7396) );
  INVX2 U8666 ( .A(length2[1]), .Y(n7423) );
  INVX2 U8667 ( .A(reg_length2[1]), .Y(n7625) );
  INVX2 U8668 ( .A(reg_length2[2]), .Y(n7626) );
  NOR4X1 U8669 ( .A(reg_length11[1]), .B(n2404), .C(n800), .D(N7871), .Y(n2472) );
  INVX2 U8670 ( .A(length4[1]), .Y(n7404) );
  INVX2 U8671 ( .A(length6[1]), .Y(n7390) );
  INVX2 U8672 ( .A(y_out_sum7[24]), .Y(n6869) );
  INVX2 U8673 ( .A(y_out_sum10[24]), .Y(n6971) );
  INVX2 U8674 ( .A(y_out_sum7[20]), .Y(n6872) );
  INVX2 U8675 ( .A(y_out_sum10[20]), .Y(n6974) );
  INVX2 U8676 ( .A(y_out_sum13[24]), .Y(n6821) );
  INVX2 U8677 ( .A(y_out_sum7[25]), .Y(n6870) );
  INVX2 U8678 ( .A(n724), .Y(n7256) );
  AOI22X1 U8679 ( .A0(reg_length10[3]), .A1(n725), .B0(reg_length10[2]), .B1(
        n726), .Y(n724) );
  INVX2 U8680 ( .A(y_out_sum10[25]), .Y(n6972) );
  INVX2 U8681 ( .A(y_out_sum13[20]), .Y(n6824) );
  INVX2 U8682 ( .A(y_out_sum9[24]), .Y(n6845) );
  AOI22X1 U8683 ( .A0(n7030), .A1(n2636), .B0(temp_w_mat_idx[0]), .B1(n2590), 
        .Y(n2632) );
  NAND2BX1 U8684 ( .AN(n2637), .B(n2638), .Y(n2636) );
  INVX2 U8685 ( .A(y_out_sum13[25]), .Y(n6822) );
  INVX2 U8686 ( .A(y_out_sum9[20]), .Y(n6848) );
  INVX2 U8687 ( .A(y_out_sum7[21]), .Y(n6873) );
  INVX2 U8688 ( .A(y_out_sum10[21]), .Y(n6976) );
  INVX2 U8689 ( .A(y_out_sum9[25]), .Y(n6846) );
  INVX2 U8690 ( .A(y_out_sum12[24]), .Y(n6797) );
  INVX2 U8691 ( .A(y_out_sum10[28]), .Y(n6968) );
  INVX2 U8692 ( .A(y_out_sum7[28]), .Y(n6866) );
  NOR4X1 U8693 ( .A(reg_length6[1]), .B(n2518), .C(n884), .D(N7688), .Y(n2508)
         );
  NOR4X1 U8694 ( .A(n2519), .B(reg_length06[3]), .C(reg_length06[5]), .D(
        reg_length06[4]), .Y(n2518) );
  NAND3X1 U8695 ( .A(n4948), .B(n4896), .C(reg_length06[0]), .Y(n2519) );
  INVX2 U8696 ( .A(y_out_sum13[21]), .Y(n6825) );
  INVX2 U8697 ( .A(y_out_sum12[20]), .Y(n6800) );
  INVX2 U8698 ( .A(y_out_sum13[28]), .Y(n6818) );
  INVX2 U8699 ( .A(reg_length0[0]), .Y(N7429) );
  INVX2 U8700 ( .A(y_out_sum7[29]), .Y(n6867) );
  INVX2 U8701 ( .A(y_out_sum12[25]), .Y(n6798) );
  INVX2 U8702 ( .A(reg_length6[2]), .Y(n7605) );
  INVX2 U8703 ( .A(y_out_sum9[21]), .Y(n6849) );
  INVX2 U8704 ( .A(y_out_sum9[28]), .Y(n6842) );
  INVX2 U8705 ( .A(y_out_sum10[29]), .Y(n6969) );
  INVX2 U8706 ( .A(reg_length6[1]), .Y(n7604) );
  INVX2 U8707 ( .A(y_out_sum12[21]), .Y(n6801) );
  INVX2 U8708 ( .A(y_out_sum13[29]), .Y(n6819) );
  INVX2 U8709 ( .A(y_out_sum12[28]), .Y(n6794) );
  INVX2 U8710 ( .A(y_out_sum9[29]), .Y(n6843) );
  INVX2 U8711 ( .A(n5650), .Y(n3007) );
  AOI222XL U8712 ( .A0(store_matrix7[11]), .A1(n5466), .B0(w_in3[11]), .B1(
        n5413), .C0(store_matrix3[11]), .C1(n5462), .Y(n5650) );
  INVX2 U8713 ( .A(n5651), .Y(n3006) );
  AOI222XL U8714 ( .A0(store_matrix7[12]), .A1(n5466), .B0(w_in3[12]), .B1(
        n5413), .C0(store_matrix3[12]), .C1(n5462), .Y(n5651) );
  INVX2 U8715 ( .A(n5652), .Y(n3005) );
  AOI222XL U8716 ( .A0(store_matrix7[13]), .A1(n5466), .B0(w_in3[13]), .B1(
        n5413), .C0(store_matrix3[13]), .C1(n5462), .Y(n5652) );
  INVX2 U8717 ( .A(n5653), .Y(n3004) );
  AOI222XL U8718 ( .A0(store_matrix7[14]), .A1(n5466), .B0(w_in3[14]), .B1(
        n5413), .C0(store_matrix3[14]), .C1(n5462), .Y(n5653) );
  INVX2 U8719 ( .A(n5654), .Y(n3003) );
  AOI222XL U8720 ( .A0(store_matrix7[15]), .A1(n5466), .B0(w_in3[15]), .B1(
        n5413), .C0(store_matrix3[15]), .C1(n5462), .Y(n5654) );
  INVX2 U8721 ( .A(n5655), .Y(n3082) );
  AOI222XL U8722 ( .A0(store_matrix6[0]), .A1(n5466), .B0(w_in2[0]), .B1(n5413), .C0(store_matrix2[0]), .C1(n5462), .Y(n5655) );
  INVX2 U8723 ( .A(n5656), .Y(n3081) );
  AOI222XL U8724 ( .A0(store_matrix6[1]), .A1(n5466), .B0(w_in2[1]), .B1(n5413), .C0(store_matrix2[1]), .C1(n5462), .Y(n5656) );
  INVX2 U8725 ( .A(n5657), .Y(n3080) );
  AOI222XL U8726 ( .A0(store_matrix6[2]), .A1(n5466), .B0(w_in2[2]), .B1(n5413), .C0(store_matrix2[2]), .C1(n5461), .Y(n5657) );
  INVX2 U8727 ( .A(n5658), .Y(n3079) );
  AOI222XL U8728 ( .A0(store_matrix6[3]), .A1(n5466), .B0(w_in2[3]), .B1(n5413), .C0(store_matrix2[3]), .C1(n5461), .Y(n5658) );
  INVX2 U8729 ( .A(n5659), .Y(n3078) );
  AOI222XL U8730 ( .A0(store_matrix6[4]), .A1(n5466), .B0(w_in2[4]), .B1(n5413), .C0(store_matrix2[4]), .C1(n5461), .Y(n5659) );
  INVX2 U8731 ( .A(n5660), .Y(n3077) );
  AOI222XL U8732 ( .A0(store_matrix6[5]), .A1(n5466), .B0(w_in2[5]), .B1(n5413), .C0(store_matrix2[5]), .C1(n5461), .Y(n5660) );
  INVX2 U8733 ( .A(n5663), .Y(n3074) );
  AOI222XL U8734 ( .A0(store_matrix6[8]), .A1(n5466), .B0(w_in2[8]), .B1(n5411), .C0(store_matrix2[8]), .C1(n5461), .Y(n5663) );
  INVX2 U8735 ( .A(n5664), .Y(n3073) );
  AOI222XL U8736 ( .A0(store_matrix6[9]), .A1(n5466), .B0(w_in2[9]), .B1(n5410), .C0(store_matrix2[9]), .C1(n5461), .Y(n5664) );
  INVX2 U8737 ( .A(n5665), .Y(n3072) );
  AOI222XL U8738 ( .A0(store_matrix6[10]), .A1(n5466), .B0(w_in2[10]), .B1(
        n5409), .C0(store_matrix2[10]), .C1(n5461), .Y(n5665) );
  INVX2 U8739 ( .A(n5666), .Y(n3071) );
  AOI222XL U8740 ( .A0(store_matrix6[11]), .A1(n5466), .B0(w_in2[11]), .B1(
        n5408), .C0(store_matrix2[11]), .C1(n5461), .Y(n5666) );
  INVX2 U8741 ( .A(n5667), .Y(n3070) );
  AOI222XL U8742 ( .A0(store_matrix6[12]), .A1(n5466), .B0(w_in2[12]), .B1(
        n5407), .C0(store_matrix2[12]), .C1(n5461), .Y(n5667) );
  INVX2 U8743 ( .A(n5668), .Y(n3069) );
  AOI222XL U8744 ( .A0(store_matrix6[13]), .A1(n5466), .B0(w_in2[13]), .B1(
        n5406), .C0(store_matrix2[13]), .C1(n5461), .Y(n5668) );
  INVX2 U8745 ( .A(n5669), .Y(n3068) );
  AOI222XL U8746 ( .A0(store_matrix6[14]), .A1(n5466), .B0(w_in2[14]), .B1(
        n5405), .C0(store_matrix2[14]), .C1(n5461), .Y(n5669) );
  INVX2 U8747 ( .A(n5648), .Y(n3009) );
  AOI222XL U8748 ( .A0(store_matrix7[9]), .A1(n5466), .B0(w_in3[9]), .B1(n5411), .C0(store_matrix3[9]), .C1(n5462), .Y(n5648) );
  INVX2 U8749 ( .A(n5670), .Y(n3067) );
  AOI222XL U8750 ( .A0(store_matrix6[15]), .A1(n5466), .B0(w_in2[15]), .B1(
        n5405), .C0(store_matrix2[15]), .C1(n5458), .Y(n5670) );
  INVX2 U8751 ( .A(n5661), .Y(n3076) );
  AOI222XL U8752 ( .A0(store_matrix6[6]), .A1(n5466), .B0(w_in2[6]), .B1(n5412), .C0(store_matrix2[6]), .C1(n5461), .Y(n5661) );
  INVX2 U8753 ( .A(n5662), .Y(n3075) );
  AOI222XL U8754 ( .A0(store_matrix6[7]), .A1(n5466), .B0(w_in2[7]), .B1(n5412), .C0(store_matrix2[7]), .C1(n5461), .Y(n5662) );
  INVX2 U8755 ( .A(n5639), .Y(n3018) );
  AOI222XL U8756 ( .A0(store_matrix7[0]), .A1(n5466), .B0(w_in3[0]), .B1(n5411), .C0(store_matrix3[0]), .C1(n5463), .Y(n5639) );
  INVX2 U8757 ( .A(n5649), .Y(n3008) );
  AOI222XL U8758 ( .A0(store_matrix7[10]), .A1(n5466), .B0(w_in3[10]), .B1(
        n5414), .C0(store_matrix3[10]), .C1(n5462), .Y(n5649) );
  INVX2 U8759 ( .A(n5644), .Y(n3013) );
  AOI222XL U8760 ( .A0(store_matrix7[5]), .A1(n5466), .B0(w_in3[5]), .B1(n5414), .C0(store_matrix3[5]), .C1(n5462), .Y(n5644) );
  INVX2 U8761 ( .A(n5645), .Y(n3012) );
  AOI222XL U8762 ( .A0(store_matrix7[6]), .A1(n5466), .B0(w_in3[6]), .B1(n5414), .C0(store_matrix3[6]), .C1(n5462), .Y(n5645) );
  INVX2 U8763 ( .A(n5646), .Y(n3011) );
  AOI222XL U8764 ( .A0(store_matrix7[7]), .A1(n5466), .B0(w_in3[7]), .B1(n5414), .C0(store_matrix3[7]), .C1(n5462), .Y(n5646) );
  INVX2 U8765 ( .A(n5647), .Y(n3010) );
  AOI222XL U8766 ( .A0(store_matrix7[8]), .A1(n5466), .B0(w_in3[8]), .B1(n5414), .C0(store_matrix3[8]), .C1(n5462), .Y(n5647) );
  INVX2 U8767 ( .A(n5640), .Y(n3017) );
  AOI222XL U8768 ( .A0(store_matrix7[1]), .A1(n5466), .B0(w_in3[1]), .B1(n5414), .C0(store_matrix3[1]), .C1(n5463), .Y(n5640) );
  INVX2 U8769 ( .A(n5641), .Y(n3016) );
  AOI222XL U8770 ( .A0(store_matrix7[2]), .A1(n5466), .B0(w_in3[2]), .B1(n5414), .C0(store_matrix3[2]), .C1(n5463), .Y(n5641) );
  INVX2 U8771 ( .A(n5642), .Y(n3015) );
  AOI222XL U8772 ( .A0(store_matrix7[3]), .A1(n5466), .B0(w_in3[3]), .B1(n5414), .C0(store_matrix3[3]), .C1(n5463), .Y(n5642) );
  INVX2 U8773 ( .A(n5643), .Y(n3014) );
  AOI222XL U8774 ( .A0(store_matrix7[4]), .A1(n5466), .B0(w_in3[4]), .B1(n5414), .C0(store_matrix3[4]), .C1(n5463), .Y(n5643) );
  INVX2 U8775 ( .A(y_out_sum12[29]), .Y(n6795) );
  AND4X2 U8776 ( .A(n2493), .B(reg_length0[0]), .C(n6788), .D(n7291), .Y(n2485) );
  INVX2 U8777 ( .A(y_out_sum11[36]), .Y(n6935) );
  INVX2 U8778 ( .A(y_out_sum11[37]), .Y(n6937) );
  INVX2 U8779 ( .A(y_out_sum14[32]), .Y(n6959) );
  AND4X2 U8780 ( .A(n7408), .B(n7409), .C(n2819), .D(n2491), .Y(n2414) );
  NOR3X1 U8781 ( .A(reg_length04[3]), .B(reg_length04[5]), .C(reg_length04[4]), 
        .Y(n2491) );
  INVX2 U8782 ( .A(y_out_sum11[32]), .Y(n6929) );
  INVX2 U8783 ( .A(y_out_sum14[36]), .Y(n6953) );
  NOR3X1 U8784 ( .A(reg_length8[3]), .B(reg_length8[5]), .C(reg_length8[4]), 
        .Y(n797) );
  INVX2 U8785 ( .A(y_out_sum11[33]), .Y(n6930) );
  INVX2 U8786 ( .A(y_out_sum14[33]), .Y(n6961) );
  INVX2 U8787 ( .A(y_out_sum14[37]), .Y(n6954) );
  OAI2BB2X1 U8788 ( .B0(n2858), .B1(n2365), .A0N(n2858), .A1N(n5350), .Y(n4002) );
  AOI22X1 U8789 ( .A0(reg_length14[4]), .A1(n344), .B0(reg_length10[5]), .B1(
        n345), .Y(n276) );
  OAI221X1 U8790 ( .A0(n111), .A1(n5674), .B0(n5415), .B1(n5673), .C0(n5672), 
        .Y(n3034) );
  AOI2BB2X1 U8791 ( .B0(store_matrix1[0]), .B1(n5445), .A0N(n5398), .A1N(n5671), .Y(n5672) );
  CLKINVXL U8792 ( .A(w_in1[0]), .Y(n5671) );
  OAI221X1 U8793 ( .A0(n5464), .A1(n5690), .B0(n5415), .B1(n5689), .C0(n5688), 
        .Y(n3030) );
  AOI2BB2X1 U8794 ( .B0(store_matrix1[4]), .B1(n5451), .A0N(n5399), .A1N(n5687), .Y(n5688) );
  CLKINVXL U8795 ( .A(w_in1[4]), .Y(n5687) );
  OAI221X1 U8796 ( .A0(n5464), .A1(n5694), .B0(n5415), .B1(n5693), .C0(n5692), 
        .Y(n3029) );
  AOI2BB2X1 U8797 ( .B0(store_matrix1[5]), .B1(n5452), .A0N(n5399), .A1N(n5691), .Y(n5692) );
  CLKINVXL U8798 ( .A(w_in1[5]), .Y(n5691) );
  OAI221X1 U8799 ( .A0(n5464), .A1(n5698), .B0(n5415), .B1(n5697), .C0(n5696), 
        .Y(n3028) );
  AOI2BB2X1 U8800 ( .B0(store_matrix1[6]), .B1(n5443), .A0N(n5399), .A1N(n5695), .Y(n5696) );
  CLKINVXL U8801 ( .A(w_in1[6]), .Y(n5695) );
  OAI221X1 U8802 ( .A0(n5464), .A1(n5702), .B0(n5415), .B1(n5701), .C0(n5700), 
        .Y(n3027) );
  AOI2BB2X1 U8803 ( .B0(store_matrix1[7]), .B1(n5452), .A0N(n5399), .A1N(n5699), .Y(n5700) );
  CLKINVXL U8804 ( .A(w_in1[7]), .Y(n5699) );
  OAI221X1 U8805 ( .A0(n5464), .A1(n5706), .B0(n5415), .B1(n5705), .C0(n5704), 
        .Y(n3026) );
  AOI2BB2X1 U8806 ( .B0(store_matrix1[8]), .B1(n5452), .A0N(n5399), .A1N(n5703), .Y(n5704) );
  CLKINVXL U8807 ( .A(w_in1[8]), .Y(n5703) );
  OAI221X1 U8808 ( .A0(n5464), .A1(n5710), .B0(n5415), .B1(n5709), .C0(n5708), 
        .Y(n3025) );
  AOI2BB2X1 U8809 ( .B0(store_matrix1[9]), .B1(n5444), .A0N(n5399), .A1N(n5707), .Y(n5708) );
  CLKINVXL U8810 ( .A(w_in1[9]), .Y(n5707) );
  OAI221X1 U8811 ( .A0(n5464), .A1(n5714), .B0(n5415), .B1(n5713), .C0(n5712), 
        .Y(n3024) );
  AOI2BB2X1 U8812 ( .B0(store_matrix1[10]), .B1(n5452), .A0N(n5399), .A1N(
        n5711), .Y(n5712) );
  CLKINVXL U8813 ( .A(w_in1[10]), .Y(n5711) );
  OAI221X1 U8814 ( .A0(n5464), .A1(n5718), .B0(n5415), .B1(n5717), .C0(n5716), 
        .Y(n3023) );
  AOI2BB2X1 U8815 ( .B0(store_matrix1[11]), .B1(n5452), .A0N(n5399), .A1N(
        n5715), .Y(n5716) );
  CLKINVXL U8816 ( .A(w_in1[11]), .Y(n5715) );
  OAI221X1 U8817 ( .A0(n5464), .A1(n5722), .B0(n5415), .B1(n5721), .C0(n5720), 
        .Y(n3022) );
  AOI2BB2X1 U8818 ( .B0(store_matrix1[12]), .B1(n5446), .A0N(n5399), .A1N(
        n5719), .Y(n5720) );
  CLKINVXL U8819 ( .A(w_in1[12]), .Y(n5719) );
  OAI221X1 U8820 ( .A0(n111), .A1(n5726), .B0(n5415), .B1(n5725), .C0(n5724), 
        .Y(n3021) );
  AOI2BB2X1 U8821 ( .B0(store_matrix1[13]), .B1(n5445), .A0N(n5399), .A1N(
        n5723), .Y(n5724) );
  CLKINVXL U8822 ( .A(w_in1[13]), .Y(n5723) );
  OAI221X1 U8823 ( .A0(n111), .A1(n5730), .B0(n5415), .B1(n5729), .C0(n5728), 
        .Y(n3020) );
  AOI2BB2X1 U8824 ( .B0(store_matrix1[14]), .B1(n5443), .A0N(n5399), .A1N(
        n5727), .Y(n5728) );
  CLKINVXL U8825 ( .A(w_in1[14]), .Y(n5727) );
  OAI221X1 U8826 ( .A0(n111), .A1(n5734), .B0(n5415), .B1(n5733), .C0(n5732), 
        .Y(n3019) );
  AOI2BB2X1 U8827 ( .B0(store_matrix1[15]), .B1(n5447), .A0N(n5399), .A1N(
        n5731), .Y(n5732) );
  CLKINVXL U8828 ( .A(w_in1[15]), .Y(n5731) );
  OAI221X1 U8829 ( .A0(n111), .A1(n5738), .B0(n5415), .B1(n5737), .C0(n5736), 
        .Y(n3050) );
  AOI2BB2X1 U8830 ( .B0(store_matrix0[0]), .B1(n5452), .A0N(n5399), .A1N(n5735), .Y(n5736) );
  CLKINVXL U8831 ( .A(w_in0[0]), .Y(n5735) );
  OAI221X1 U8832 ( .A0(n5464), .A1(n5686), .B0(n5415), .B1(n5685), .C0(n5684), 
        .Y(n3031) );
  AOI2BB2X1 U8833 ( .B0(store_matrix1[3]), .B1(n5446), .A0N(n5399), .A1N(n5683), .Y(n5684) );
  CLKINVXL U8834 ( .A(w_in1[3]), .Y(n5683) );
  OAI221X1 U8835 ( .A0(n111), .A1(n5742), .B0(n5415), .B1(n5741), .C0(n5740), 
        .Y(n3049) );
  AOI2BB2X1 U8836 ( .B0(store_matrix0[1]), .B1(n5453), .A0N(n5399), .A1N(n5739), .Y(n5740) );
  CLKINVXL U8837 ( .A(w_in0[1]), .Y(n5739) );
  OAI221X1 U8838 ( .A0(n111), .A1(n5746), .B0(n5415), .B1(n5745), .C0(n5744), 
        .Y(n3048) );
  AOI2BB2X1 U8839 ( .B0(store_matrix0[2]), .B1(n5448), .A0N(n5399), .A1N(n5743), .Y(n5744) );
  CLKINVXL U8840 ( .A(w_in0[2]), .Y(n5743) );
  OAI221X1 U8841 ( .A0(n111), .A1(n5750), .B0(n5415), .B1(n5749), .C0(n5748), 
        .Y(n3047) );
  AOI2BB2X1 U8842 ( .B0(store_matrix0[3]), .B1(n5453), .A0N(n5399), .A1N(n5747), .Y(n5748) );
  CLKINVXL U8843 ( .A(w_in0[3]), .Y(n5747) );
  OAI221X1 U8844 ( .A0(n111), .A1(n5754), .B0(n5415), .B1(n5753), .C0(n5752), 
        .Y(n3046) );
  AOI2BB2X1 U8845 ( .B0(store_matrix0[4]), .B1(n5447), .A0N(n5399), .A1N(n5751), .Y(n5752) );
  CLKINVXL U8846 ( .A(w_in0[4]), .Y(n5751) );
  OAI221X1 U8847 ( .A0(n111), .A1(n5758), .B0(n5415), .B1(n5757), .C0(n5756), 
        .Y(n3045) );
  AOI2BB2X1 U8848 ( .B0(store_matrix0[5]), .B1(n5449), .A0N(n5399), .A1N(n5755), .Y(n5756) );
  CLKINVXL U8849 ( .A(w_in0[5]), .Y(n5755) );
  OAI221X1 U8850 ( .A0(n111), .A1(n5762), .B0(n5415), .B1(n5761), .C0(n5760), 
        .Y(n3044) );
  AOI2BB2X1 U8851 ( .B0(store_matrix0[6]), .B1(n5454), .A0N(n5399), .A1N(n5759), .Y(n5760) );
  CLKINVXL U8852 ( .A(w_in0[6]), .Y(n5759) );
  OAI221X1 U8853 ( .A0(n111), .A1(n5766), .B0(n5415), .B1(n5765), .C0(n5764), 
        .Y(n3043) );
  AOI2BB2X1 U8854 ( .B0(store_matrix0[7]), .B1(n5454), .A0N(n5399), .A1N(n5763), .Y(n5764) );
  CLKINVXL U8855 ( .A(w_in0[7]), .Y(n5763) );
  OAI221X1 U8856 ( .A0(n111), .A1(n5770), .B0(n5415), .B1(n5769), .C0(n5768), 
        .Y(n3042) );
  AOI2BB2X1 U8857 ( .B0(store_matrix0[8]), .B1(n5449), .A0N(n5399), .A1N(n5767), .Y(n5768) );
  CLKINVXL U8858 ( .A(w_in0[8]), .Y(n5767) );
  OAI221X1 U8859 ( .A0(n111), .A1(n5774), .B0(n5415), .B1(n5773), .C0(n5772), 
        .Y(n3041) );
  AOI2BB2X1 U8860 ( .B0(store_matrix0[9]), .B1(n5455), .A0N(n5399), .A1N(n5771), .Y(n5772) );
  CLKINVXL U8861 ( .A(w_in0[9]), .Y(n5771) );
  OAI221X1 U8862 ( .A0(n111), .A1(n5778), .B0(n5415), .B1(n5777), .C0(n5776), 
        .Y(n3040) );
  AOI2BB2X1 U8863 ( .B0(store_matrix0[10]), .B1(n5455), .A0N(n5399), .A1N(
        n5775), .Y(n5776) );
  CLKINVXL U8864 ( .A(w_in0[10]), .Y(n5775) );
  OAI221X1 U8865 ( .A0(n111), .A1(n5782), .B0(n5415), .B1(n5781), .C0(n5780), 
        .Y(n3039) );
  AOI2BB2X1 U8866 ( .B0(store_matrix0[11]), .B1(n5444), .A0N(n5399), .A1N(
        n5779), .Y(n5780) );
  CLKINVXL U8867 ( .A(w_in0[11]), .Y(n5779) );
  OAI221X1 U8868 ( .A0(n111), .A1(n5786), .B0(n5415), .B1(n5785), .C0(n5784), 
        .Y(n3038) );
  AOI2BB2X1 U8869 ( .B0(store_matrix0[12]), .B1(n5456), .A0N(n5399), .A1N(
        n5783), .Y(n5784) );
  CLKINVXL U8870 ( .A(w_in0[12]), .Y(n5783) );
  OAI221X1 U8871 ( .A0(n111), .A1(n5790), .B0(n5415), .B1(n5789), .C0(n5788), 
        .Y(n3037) );
  AOI2BB2X1 U8872 ( .B0(store_matrix0[13]), .B1(n5456), .A0N(n5399), .A1N(
        n5787), .Y(n5788) );
  CLKINVXL U8873 ( .A(w_in0[13]), .Y(n5787) );
  OAI221X1 U8874 ( .A0(n111), .A1(n5794), .B0(n5415), .B1(n5793), .C0(n5792), 
        .Y(n3036) );
  AOI2BB2X1 U8875 ( .B0(store_matrix0[14]), .B1(n5450), .A0N(n5399), .A1N(
        n5791), .Y(n5792) );
  CLKINVXL U8876 ( .A(w_in0[14]), .Y(n5791) );
  OAI221X1 U8877 ( .A0(n111), .A1(n5798), .B0(n5415), .B1(n5797), .C0(n5796), 
        .Y(n3035) );
  AOI2BB2X1 U8878 ( .B0(store_matrix0[15]), .B1(n5448), .A0N(n5399), .A1N(
        n5795), .Y(n5796) );
  CLKINVXL U8879 ( .A(w_in0[15]), .Y(n5795) );
  OAI221X1 U8880 ( .A0(n5464), .A1(n5678), .B0(n5415), .B1(n5677), .C0(n5676), 
        .Y(n3033) );
  AOI2BB2X1 U8881 ( .B0(store_matrix1[1]), .B1(n5450), .A0N(n5400), .A1N(n5675), .Y(n5676) );
  CLKINVXL U8882 ( .A(w_in1[1]), .Y(n5675) );
  OAI221X1 U8883 ( .A0(n5464), .A1(n5682), .B0(n5415), .B1(n5681), .C0(n5680), 
        .Y(n3032) );
  AOI2BB2X1 U8884 ( .B0(store_matrix1[2]), .B1(n5451), .A0N(n5400), .A1N(n5679), .Y(n5680) );
  CLKINVXL U8885 ( .A(w_in1[2]), .Y(n5679) );
  NOR3X1 U8886 ( .A(reg_length11[3]), .B(reg_length11[5]), .C(reg_length11[4]), 
        .Y(n799) );
  NOR3X1 U8887 ( .A(reg_length7[3]), .B(reg_length7[5]), .C(reg_length7[4]), 
        .Y(n849) );
  AND4X2 U8888 ( .A(n7436), .B(n7437), .C(n2816), .D(n2506), .Y(n2420) );
  NOR3X1 U8889 ( .A(reg_length01[3]), .B(reg_length01[5]), .C(reg_length01[4]), 
        .Y(n2506) );
  NAND4X1 U8890 ( .A(n7400), .B(n7401), .C(n2820), .D(n2504), .Y(n2417) );
  NOR3X1 U8891 ( .A(reg_length05[3]), .B(reg_length05[5]), .C(reg_length05[4]), 
        .Y(n2504) );
  OAI2BB1X1 U8892 ( .A0N(Q32[13]), .A1N(n5349), .B0(n5876), .Y(n2910) );
  OAI2BB1X1 U8893 ( .A0N(Q42[10]), .A1N(n5445), .B0(n5857), .Y(n2929) );
  OAI2BB1X1 U8894 ( .A0N(Q42[11]), .A1N(n5444), .B0(n5858), .Y(n2928) );
  OAI2BB1X1 U8895 ( .A0N(Q42[12]), .A1N(n5459), .B0(n5859), .Y(n2927) );
  OAI2BB1X1 U8896 ( .A0N(Q42[13]), .A1N(n5443), .B0(n5860), .Y(n2926) );
  OAI2BB1X1 U8897 ( .A0N(Q42[14]), .A1N(n5456), .B0(n5861), .Y(n2925) );
  OAI2BB1X1 U8898 ( .A0N(Q42[1]), .A1N(n5449), .B0(n5848), .Y(n2938) );
  OAI2BB1X1 U8899 ( .A0N(Q42[2]), .A1N(n5448), .B0(n5849), .Y(n2937) );
  OAI2BB1X1 U8900 ( .A0N(Q42[3]), .A1N(n5460), .B0(n5850), .Y(n2936) );
  OAI2BB1X1 U8901 ( .A0N(Q42[4]), .A1N(n5447), .B0(n5851), .Y(n2935) );
  OAI2BB1X1 U8902 ( .A0N(Q42[5]), .A1N(n5460), .B0(n5852), .Y(n2934) );
  OAI2BB1X1 U8903 ( .A0N(Q42[6]), .A1N(n5459), .B0(n5853), .Y(n2933) );
  OAI2BB1X1 U8904 ( .A0N(Q42[7]), .A1N(n5460), .B0(n5854), .Y(n2932) );
  OAI2BB1X1 U8905 ( .A0N(Q42[8]), .A1N(n5446), .B0(n5855), .Y(n2931) );
  OAI2BB1X1 U8906 ( .A0N(Q42[9]), .A1N(n5459), .B0(n5856), .Y(n2930) );
  OAI2BB1X1 U8907 ( .A0N(Q62[11]), .A1N(n5460), .B0(n5826), .Y(n2960) );
  OAI2BB1X1 U8908 ( .A0N(Q62[12]), .A1N(n5460), .B0(n5827), .Y(n2959) );
  OAI2BB1X1 U8909 ( .A0N(Q62[13]), .A1N(n5460), .B0(n5828), .Y(n2958) );
  OAI2BB1X1 U8910 ( .A0N(Q62[14]), .A1N(n5460), .B0(n5829), .Y(n2957) );
  OAI2BB1X1 U8911 ( .A0N(Q62[15]), .A1N(n5460), .B0(n5830), .Y(n2956) );
  OAI2BB1X1 U8912 ( .A0N(Q52[10]), .A1N(n5460), .B0(n5841), .Y(n2945) );
  OAI2BB1X1 U8913 ( .A0N(Q52[11]), .A1N(n5452), .B0(n5842), .Y(n2944) );
  OAI2BB1X1 U8914 ( .A0N(Q52[12]), .A1N(n5452), .B0(n5843), .Y(n2943) );
  OAI2BB1X1 U8915 ( .A0N(Q52[13]), .A1N(n5460), .B0(n5844), .Y(n2942) );
  OAI2BB1X1 U8916 ( .A0N(Q52[14]), .A1N(n5451), .B0(n5845), .Y(n2941) );
  OAI2BB1X1 U8917 ( .A0N(Q52[15]), .A1N(n5450), .B0(n5846), .Y(n2940) );
  OAI2BB1X1 U8918 ( .A0N(Q52[1]), .A1N(n5460), .B0(n5832), .Y(n2954) );
  OAI2BB1X1 U8919 ( .A0N(Q52[2]), .A1N(n5460), .B0(n5833), .Y(n2953) );
  OAI2BB1X1 U8920 ( .A0N(Q52[3]), .A1N(n5455), .B0(n5834), .Y(n2952) );
  OAI2BB1X1 U8921 ( .A0N(Q52[4]), .A1N(n5460), .B0(n5835), .Y(n2951) );
  OAI2BB1X1 U8922 ( .A0N(Q52[5]), .A1N(n5454), .B0(n5836), .Y(n2950) );
  OAI2BB1X1 U8923 ( .A0N(Q52[6]), .A1N(n5453), .B0(n5837), .Y(n2949) );
  OAI2BB1X1 U8924 ( .A0N(Q52[7]), .A1N(n5460), .B0(n5838), .Y(n2948) );
  OAI2BB1X1 U8925 ( .A0N(Q52[8]), .A1N(n5452), .B0(n5839), .Y(n2947) );
  OAI2BB1X1 U8926 ( .A0N(Q52[9]), .A1N(n5460), .B0(n5840), .Y(n2946) );
  OAI2BB1X1 U8927 ( .A0N(Q42[0]), .A1N(n5460), .B0(n5847), .Y(n2939) );
  OR2X1 U8928 ( .A(n5401), .B(n5471), .Y(n5847) );
  OAI2BB1X1 U8929 ( .A0N(Q52[0]), .A1N(n5460), .B0(n5831), .Y(n2955) );
  OR2X1 U8930 ( .A(n5401), .B(n5470), .Y(n5831) );
  OAI2BB1X1 U8931 ( .A0N(Q22[10]), .A1N(n5895), .B0(n5889), .Y(n2897) );
  OAI2BB1X1 U8932 ( .A0N(Q22[11]), .A1N(n5348), .B0(n5890), .Y(n2896) );
  OAI2BB1X1 U8933 ( .A0N(Q22[12]), .A1N(n5349), .B0(n5891), .Y(n2895) );
  OAI2BB1X1 U8934 ( .A0N(Q22[13]), .A1N(n5895), .B0(n5892), .Y(n2894) );
  OAI2BB1X1 U8935 ( .A0N(Q22[14]), .A1N(n5348), .B0(n5893), .Y(n2893) );
  OAI2BB1X1 U8936 ( .A0N(Q22[15]), .A1N(n5349), .B0(n5894), .Y(n2892) );
  OAI2BB1X1 U8937 ( .A0N(Q22[1]), .A1N(n5895), .B0(n5880), .Y(n2906) );
  OAI2BB1X1 U8938 ( .A0N(Q22[2]), .A1N(n5348), .B0(n5881), .Y(n2905) );
  OAI2BB1X1 U8939 ( .A0N(Q22[3]), .A1N(n5349), .B0(n5882), .Y(n2904) );
  OAI2BB1X1 U8940 ( .A0N(Q22[4]), .A1N(n5895), .B0(n5883), .Y(n2903) );
  OAI2BB1X1 U8941 ( .A0N(Q22[5]), .A1N(n5348), .B0(n5884), .Y(n2902) );
  OAI2BB1X1 U8942 ( .A0N(Q22[6]), .A1N(n5349), .B0(n5885), .Y(n2901) );
  OAI2BB1X1 U8943 ( .A0N(Q22[7]), .A1N(n5895), .B0(n5886), .Y(n2900) );
  OAI2BB1X1 U8944 ( .A0N(Q22[8]), .A1N(n5348), .B0(n5887), .Y(n2899) );
  OAI2BB1X1 U8945 ( .A0N(Q22[9]), .A1N(n5349), .B0(n5888), .Y(n2898) );
  OAI2BB1X1 U8946 ( .A0N(Q32[10]), .A1N(n5349), .B0(n5873), .Y(n2913) );
  OAI2BB1X1 U8947 ( .A0N(Q32[11]), .A1N(n5895), .B0(n5874), .Y(n2912) );
  OAI2BB1X1 U8948 ( .A0N(Q32[12]), .A1N(n5348), .B0(n5875), .Y(n2911) );
  OAI2BB1X1 U8949 ( .A0N(Q32[14]), .A1N(n5895), .B0(n5877), .Y(n2909) );
  OAI2BB1X1 U8950 ( .A0N(Q32[15]), .A1N(n5348), .B0(n5878), .Y(n2908) );
  OAI2BB1X1 U8951 ( .A0N(Q32[1]), .A1N(n5349), .B0(n5864), .Y(n2922) );
  OAI2BB1X1 U8952 ( .A0N(Q32[2]), .A1N(n5895), .B0(n5865), .Y(n2921) );
  OAI2BB1X1 U8953 ( .A0N(Q32[3]), .A1N(n5348), .B0(n5866), .Y(n2920) );
  OAI2BB1X1 U8954 ( .A0N(Q32[4]), .A1N(n5349), .B0(n5867), .Y(n2919) );
  OAI2BB1X1 U8955 ( .A0N(Q32[5]), .A1N(n5895), .B0(n5868), .Y(n2918) );
  OAI2BB1X1 U8956 ( .A0N(Q32[6]), .A1N(n5348), .B0(n5869), .Y(n2917) );
  OAI2BB1X1 U8957 ( .A0N(Q32[7]), .A1N(n5349), .B0(n5870), .Y(n2916) );
  OAI2BB1X1 U8958 ( .A0N(Q32[8]), .A1N(n5895), .B0(n5871), .Y(n2915) );
  OAI2BB1X1 U8959 ( .A0N(Q32[9]), .A1N(n5348), .B0(n5872), .Y(n2914) );
  OAI2BB1X1 U8960 ( .A0N(Q22[0]), .A1N(n5349), .B0(n5879), .Y(n2907) );
  OR2X1 U8961 ( .A(n5400), .B(n5473), .Y(n5879) );
  OAI2BB1X1 U8962 ( .A0N(Q32[0]), .A1N(n5348), .B0(n5863), .Y(n2923) );
  OR2X1 U8963 ( .A(n5400), .B(n5472), .Y(n5863) );
  OAI2BB1X1 U8964 ( .A0N(Q42[15]), .A1N(n5460), .B0(n5862), .Y(n2924) );
  OAI2BB1X1 U8965 ( .A0N(Q72[0]), .A1N(n5460), .B0(n5799), .Y(n2986) );
  OR2X1 U8966 ( .A(n5400), .B(n5468), .Y(n5799) );
  AND4X2 U8967 ( .A(n4946), .B(n4894), .C(reg_length08[0]), .D(n2492), .Y(
        n2418) );
  NOR3X1 U8968 ( .A(reg_length08[3]), .B(reg_length08[5]), .C(reg_length08[4]), 
        .Y(n2492) );
  INVX2 U8969 ( .A(y_out_sum10[32]), .Y(n6962) );
  NAND4X1 U8970 ( .A(n7428), .B(n7429), .C(n2817), .D(n2505), .Y(n2413) );
  NOR3X1 U8971 ( .A(reg_length02[3]), .B(reg_length02[5]), .C(reg_length02[4]), 
        .Y(n2505) );
  INVX2 U8972 ( .A(y_out_sum10[36]), .Y(n6965) );
  OAI2BB1X1 U8973 ( .A0N(Q62[10]), .A1N(n5460), .B0(n5825), .Y(n2961) );
  OAI2BB1X1 U8974 ( .A0N(Q62[1]), .A1N(n5460), .B0(n5816), .Y(n2970) );
  OAI2BB1X1 U8975 ( .A0N(Q62[2]), .A1N(n5460), .B0(n5817), .Y(n2969) );
  OAI2BB1X1 U8976 ( .A0N(Q62[3]), .A1N(n5460), .B0(n5818), .Y(n2968) );
  OAI2BB1X1 U8977 ( .A0N(Q62[4]), .A1N(n5460), .B0(n5819), .Y(n2967) );
  OAI2BB1X1 U8978 ( .A0N(Q62[5]), .A1N(n5460), .B0(n5820), .Y(n2966) );
  OAI2BB1X1 U8979 ( .A0N(Q62[6]), .A1N(n5460), .B0(n5821), .Y(n2965) );
  OAI2BB1X1 U8980 ( .A0N(Q62[7]), .A1N(n5460), .B0(n5822), .Y(n2964) );
  OAI2BB1X1 U8981 ( .A0N(Q62[8]), .A1N(n5460), .B0(n5823), .Y(n2963) );
  OAI2BB1X1 U8982 ( .A0N(Q62[9]), .A1N(n5460), .B0(n5824), .Y(n2962) );
  OAI2BB1X1 U8983 ( .A0N(Q72[10]), .A1N(n5460), .B0(n5809), .Y(n2976) );
  OAI2BB1X1 U8984 ( .A0N(Q72[11]), .A1N(n5460), .B0(n5810), .Y(n2975) );
  OAI2BB1X1 U8985 ( .A0N(Q72[12]), .A1N(n5460), .B0(n5811), .Y(n2974) );
  OAI2BB1X1 U8986 ( .A0N(Q72[13]), .A1N(n5460), .B0(n5812), .Y(n2973) );
  OAI2BB1X1 U8987 ( .A0N(Q72[14]), .A1N(n5460), .B0(n5813), .Y(n2972) );
  OAI2BB1X1 U8988 ( .A0N(Q72[15]), .A1N(n5460), .B0(n5814), .Y(n2971) );
  OAI2BB1X1 U8989 ( .A0N(Q72[1]), .A1N(n5460), .B0(n5800), .Y(n2985) );
  OAI2BB1X1 U8990 ( .A0N(Q72[2]), .A1N(n5460), .B0(n5801), .Y(n2984) );
  OAI2BB1X1 U8991 ( .A0N(Q72[3]), .A1N(n5460), .B0(n5802), .Y(n2983) );
  OAI2BB1X1 U8992 ( .A0N(Q72[4]), .A1N(n5460), .B0(n5803), .Y(n2982) );
  OAI2BB1X1 U8993 ( .A0N(Q72[5]), .A1N(n5460), .B0(n5804), .Y(n2981) );
  OAI2BB1X1 U8994 ( .A0N(Q72[6]), .A1N(n5460), .B0(n5805), .Y(n2980) );
  OAI2BB1X1 U8995 ( .A0N(Q72[7]), .A1N(n5460), .B0(n5806), .Y(n2979) );
  OAI2BB1X1 U8996 ( .A0N(Q72[8]), .A1N(n5460), .B0(n5807), .Y(n2978) );
  OAI2BB1X1 U8997 ( .A0N(Q72[9]), .A1N(n5460), .B0(n5808), .Y(n2977) );
  OAI2BB1X1 U8998 ( .A0N(Q62[0]), .A1N(n5460), .B0(n5815), .Y(n4029) );
  OR2X1 U8999 ( .A(n5396), .B(n5469), .Y(n5815) );
  AOI222XL U9000 ( .A0(reg_length13[3]), .A1(n7257), .B0(reg_length13[5]), 
        .B1(n7260), .C0(reg_length13[4]), .C1(n7244), .Y(n168) );
  INVX2 U9001 ( .A(y_out_sum10[37]), .Y(n6966) );
  INVX2 U9002 ( .A(y_out_sum10[33]), .Y(n6963) );
  INVX2 U9003 ( .A(y_out_sum8[36]), .Y(n6911) );
  AND4X2 U9004 ( .A(n7416), .B(n7417), .C(n2818), .D(n2507), .Y(n2415) );
  NOR3X1 U9005 ( .A(reg_length03[3]), .B(reg_length03[5]), .C(reg_length03[4]), 
        .Y(n2507) );
  INVX2 U9006 ( .A(y_out_sum8[37]), .Y(n6913) );
  AND4X2 U9007 ( .A(n4947), .B(n4895), .C(reg_length012[0]), .D(n2483), .Y(
        n2398) );
  NOR3X1 U9008 ( .A(reg_length012[3]), .B(reg_length012[5]), .C(
        reg_length012[4]), .Y(n2483) );
  INVX2 U9009 ( .A(y_out_sum8[32]), .Y(n6905) );
  OAI33X1 U9010 ( .A0(n2273), .A1(count1[0]), .A2(n802), .B0(n2533), .B1(n2534), .B2(n2535), .Y(n2527) );
  OR2X1 U9011 ( .A(n2841), .B(n2840), .Y(n2535) );
  INVX2 U9012 ( .A(y_out_sum8[33]), .Y(n6906) );
  NAND4X1 U9013 ( .A(n4949), .B(n4897), .C(reg_length010[0]), .D(n2482), .Y(
        n2401) );
  NOR3X1 U9014 ( .A(reg_length010[3]), .B(reg_length010[5]), .C(
        reg_length010[4]), .Y(n2482) );
  NOR2X1 U9015 ( .A(n103), .B(n104), .Y(n99) );
  AOI32X1 U9016 ( .A0(n7312), .A1(n7313), .A2(n107), .B0(n108), .B1(n7315), 
        .Y(n103) );
  OAI33X1 U9017 ( .A0(n7312), .A1(count[13]), .A2(n5415), .B0(n7313), .B1(
        n5378), .B2(n5464), .Y(n108) );
  NOR2X1 U9018 ( .A(n5441), .B(n7315), .Y(n107) );
  OAI22X1 U9019 ( .A0(n5396), .A1(n5588), .B0(n5440), .B1(n5725), .Y(n7163) );
  CLKINVXL U9020 ( .A(w_in7[13]), .Y(n5588) );
  OAI22X1 U9021 ( .A0(n5396), .A1(n5589), .B0(n5440), .B1(n5729), .Y(n7162) );
  CLKINVXL U9022 ( .A(w_in7[14]), .Y(n5589) );
  OAI22X1 U9023 ( .A0(n5396), .A1(n5590), .B0(n5440), .B1(n5733), .Y(n7161) );
  CLKINVXL U9024 ( .A(w_in7[15]), .Y(n5590) );
  OAI22X1 U9025 ( .A0(n5396), .A1(n5591), .B0(n5440), .B1(n5737), .Y(n7160) );
  CLKINVXL U9026 ( .A(w_in6[0]), .Y(n5591) );
  OAI22X1 U9027 ( .A0(n5396), .A1(n5592), .B0(n5440), .B1(n5741), .Y(n7159) );
  CLKINVXL U9028 ( .A(w_in6[1]), .Y(n5592) );
  OAI22X1 U9029 ( .A0(n5396), .A1(n5593), .B0(n5440), .B1(n5745), .Y(n7158) );
  CLKINVXL U9030 ( .A(w_in6[2]), .Y(n5593) );
  OAI22X1 U9031 ( .A0(n5396), .A1(n5594), .B0(n5440), .B1(n5749), .Y(n7157) );
  CLKINVXL U9032 ( .A(w_in6[3]), .Y(n5594) );
  OAI22X1 U9033 ( .A0(n5396), .A1(n5595), .B0(n5440), .B1(n5753), .Y(n7155) );
  CLKINVXL U9034 ( .A(w_in6[4]), .Y(n5595) );
  OAI22X1 U9035 ( .A0(n5396), .A1(n5596), .B0(n5440), .B1(n5757), .Y(n7154) );
  CLKINVXL U9036 ( .A(w_in6[5]), .Y(n5596) );
  OAI22X1 U9037 ( .A0(n5396), .A1(n5597), .B0(n5440), .B1(n5761), .Y(n7153) );
  CLKINVXL U9038 ( .A(w_in6[6]), .Y(n5597) );
  OAI22X1 U9039 ( .A0(n5396), .A1(n5598), .B0(n5440), .B1(n5765), .Y(n7152) );
  OAI22X1 U9040 ( .A0(n5396), .A1(n5599), .B0(n5440), .B1(n5769), .Y(n7151) );
  CLKINVXL U9041 ( .A(w_in6[8]), .Y(n5599) );
  OAI22X1 U9042 ( .A0(n5397), .A1(n5601), .B0(n5439), .B1(n5777), .Y(n7149) );
  CLKINVXL U9043 ( .A(w_in6[10]), .Y(n5601) );
  OAI22X1 U9044 ( .A0(n5396), .A1(n5602), .B0(n5439), .B1(n5781), .Y(n7148) );
  CLKINVXL U9045 ( .A(w_in6[11]), .Y(n5602) );
  OAI22X1 U9046 ( .A0(n5397), .A1(n5603), .B0(n5439), .B1(n5785), .Y(n7147) );
  CLKINVXL U9047 ( .A(w_in6[12]), .Y(n5603) );
  OAI22X1 U9048 ( .A0(n5397), .A1(n5604), .B0(n5439), .B1(n5789), .Y(n7146) );
  CLKINVXL U9049 ( .A(w_in6[13]), .Y(n5604) );
  OAI22X1 U9050 ( .A0(n5396), .A1(n5605), .B0(n5439), .B1(n5793), .Y(n7144) );
  CLKINVXL U9051 ( .A(w_in6[14]), .Y(n5605) );
  OAI22X1 U9052 ( .A0(n5397), .A1(n5606), .B0(n5439), .B1(n5797), .Y(n7143) );
  CLKINVXL U9053 ( .A(w_in6[15]), .Y(n5606) );
  OAI22X1 U9054 ( .A0(n5397), .A1(n5607), .B0(n5439), .B1(n5674), .Y(n3098) );
  CLKINVXL U9055 ( .A(w_in5[0]), .Y(n5607) );
  OAI22X1 U9056 ( .A0(n5396), .A1(n5608), .B0(n5439), .B1(n5678), .Y(n3097) );
  CLKINVXL U9057 ( .A(w_in5[1]), .Y(n5608) );
  OAI22X1 U9058 ( .A0(n5396), .A1(n5609), .B0(n5439), .B1(n5682), .Y(n3096) );
  CLKINVXL U9059 ( .A(w_in5[2]), .Y(n5609) );
  OAI22X1 U9060 ( .A0(n5397), .A1(n5610), .B0(n5439), .B1(n5686), .Y(n3095) );
  CLKINVXL U9061 ( .A(w_in5[3]), .Y(n5610) );
  OAI22X1 U9062 ( .A0(n5396), .A1(n5611), .B0(n5439), .B1(n5690), .Y(n3094) );
  CLKINVXL U9063 ( .A(w_in5[4]), .Y(n5611) );
  OAI22X1 U9064 ( .A0(n5397), .A1(n5612), .B0(n5439), .B1(n5694), .Y(n3093) );
  CLKINVXL U9065 ( .A(w_in5[5]), .Y(n5612) );
  OAI22X1 U9066 ( .A0(n5396), .A1(n5613), .B0(n5438), .B1(n5698), .Y(n3092) );
  CLKINVXL U9067 ( .A(w_in5[6]), .Y(n5613) );
  OAI22X1 U9068 ( .A0(n5397), .A1(n5614), .B0(n5438), .B1(n5702), .Y(n3091) );
  CLKINVXL U9069 ( .A(w_in5[7]), .Y(n5614) );
  OAI22X1 U9070 ( .A0(n5397), .A1(n5615), .B0(n5438), .B1(n5706), .Y(n3090) );
  CLKINVXL U9071 ( .A(w_in5[8]), .Y(n5615) );
  OAI22X1 U9072 ( .A0(n5397), .A1(n5616), .B0(n5438), .B1(n5710), .Y(n3089) );
  CLKINVXL U9073 ( .A(w_in5[9]), .Y(n5616) );
  OAI22X1 U9074 ( .A0(n5397), .A1(n5617), .B0(n5438), .B1(n5714), .Y(n3088) );
  CLKINVXL U9075 ( .A(w_in5[10]), .Y(n5617) );
  OAI22X1 U9076 ( .A0(n5397), .A1(n5618), .B0(n5438), .B1(n5718), .Y(n3087) );
  CLKINVXL U9077 ( .A(w_in5[11]), .Y(n5618) );
  OAI22X1 U9078 ( .A0(n5397), .A1(n5619), .B0(n5438), .B1(n5722), .Y(n3086) );
  CLKINVXL U9079 ( .A(w_in5[12]), .Y(n5619) );
  OAI22X1 U9080 ( .A0(n5397), .A1(n5620), .B0(n5438), .B1(n5726), .Y(n3085) );
  CLKINVXL U9081 ( .A(w_in5[13]), .Y(n5620) );
  OAI22X1 U9082 ( .A0(n5397), .A1(n5621), .B0(n5438), .B1(n5730), .Y(n3084) );
  CLKINVXL U9083 ( .A(w_in5[14]), .Y(n5621) );
  OAI22X1 U9084 ( .A0(n5397), .A1(n5622), .B0(n5438), .B1(n5734), .Y(n3083) );
  CLKINVXL U9085 ( .A(w_in5[15]), .Y(n5622) );
  OAI22X1 U9086 ( .A0(n5397), .A1(n5623), .B0(n5438), .B1(n5738), .Y(n3114) );
  CLKINVXL U9087 ( .A(w_in4[0]), .Y(n5623) );
  OAI22X1 U9088 ( .A0(n5397), .A1(n5624), .B0(n5438), .B1(n5742), .Y(n3113) );
  CLKINVXL U9089 ( .A(w_in4[1]), .Y(n5624) );
  OAI22X1 U9090 ( .A0(n5397), .A1(n5625), .B0(n5438), .B1(n5746), .Y(n3112) );
  CLKINVXL U9091 ( .A(w_in4[2]), .Y(n5625) );
  OAI22X1 U9092 ( .A0(n5397), .A1(n5626), .B0(n5437), .B1(n5750), .Y(n3111) );
  CLKINVXL U9093 ( .A(w_in4[3]), .Y(n5626) );
  NOR3X1 U9094 ( .A(reg_length13[3]), .B(reg_length13[5]), .C(reg_length13[4]), 
        .Y(n846) );
  NAND4X1 U9095 ( .A(n4950), .B(n4898), .C(reg_length09[0]), .D(n2481), .Y(
        n2402) );
  NOR3X1 U9096 ( .A(reg_length09[3]), .B(reg_length09[5]), .C(reg_length09[4]), 
        .Y(n2481) );
  INVX2 U9097 ( .A(reg_length8[2]), .Y(n7592) );
  OAI22X1 U9098 ( .A0(n5398), .A1(n5627), .B0(n5439), .B1(n5754), .Y(n3110) );
  CLKINVXL U9099 ( .A(w_in4[4]), .Y(n5627) );
  OAI22X1 U9100 ( .A0(n5398), .A1(n5629), .B0(n5437), .B1(n5762), .Y(n3108) );
  CLKINVXL U9101 ( .A(w_in4[6]), .Y(n5629) );
  OAI22X1 U9102 ( .A0(n5398), .A1(n5631), .B0(n5437), .B1(n5770), .Y(n3106) );
  CLKINVXL U9103 ( .A(w_in4[8]), .Y(n5631) );
  OAI22X1 U9104 ( .A0(n5398), .A1(n5632), .B0(n5437), .B1(n5774), .Y(n3105) );
  CLKINVXL U9105 ( .A(w_in4[9]), .Y(n5632) );
  OAI22X1 U9106 ( .A0(n5398), .A1(n5633), .B0(n5437), .B1(n5778), .Y(n3104) );
  CLKINVXL U9107 ( .A(w_in4[10]), .Y(n5633) );
  OAI22X1 U9108 ( .A0(n5398), .A1(n5634), .B0(n5437), .B1(n5782), .Y(n3103) );
  CLKINVXL U9109 ( .A(w_in4[11]), .Y(n5634) );
  OAI22X1 U9110 ( .A0(n5398), .A1(n5635), .B0(n5437), .B1(n5786), .Y(n3102) );
  CLKINVXL U9111 ( .A(w_in4[12]), .Y(n5635) );
  OAI22X1 U9112 ( .A0(n5398), .A1(n5636), .B0(n5437), .B1(n5790), .Y(n3101) );
  CLKINVXL U9113 ( .A(w_in4[13]), .Y(n5636) );
  OAI22X1 U9114 ( .A0(n5398), .A1(n5637), .B0(n5437), .B1(n5794), .Y(n3100) );
  CLKINVXL U9115 ( .A(w_in4[14]), .Y(n5637) );
  OAI22X1 U9116 ( .A0(n5398), .A1(n5638), .B0(n5437), .B1(n5798), .Y(n3099) );
  CLKINVXL U9117 ( .A(w_in4[15]), .Y(n5638) );
  OAI22X1 U9118 ( .A0(n5396), .A1(n5575), .B0(n5437), .B1(n5673), .Y(n7167) );
  CLKINVXL U9119 ( .A(w_in7[0]), .Y(n5575) );
  OAI22X1 U9120 ( .A0(n5396), .A1(n5585), .B0(n5441), .B1(n5713), .Y(n7166) );
  CLKINVXL U9121 ( .A(w_in7[10]), .Y(n5585) );
  OAI22X1 U9122 ( .A0(n5396), .A1(n5586), .B0(n5441), .B1(n5717), .Y(n7165) );
  CLKINVXL U9123 ( .A(w_in7[11]), .Y(n5586) );
  OAI22X1 U9124 ( .A0(n5397), .A1(n5587), .B0(n5441), .B1(n5721), .Y(n7164) );
  CLKINVXL U9125 ( .A(w_in7[12]), .Y(n5587) );
  OAI22X1 U9126 ( .A0(n5397), .A1(n5577), .B0(n5441), .B1(n5681), .Y(n7145) );
  CLKINVXL U9127 ( .A(w_in7[2]), .Y(n5577) );
  OAI22X1 U9128 ( .A0(n5396), .A1(n5578), .B0(n5441), .B1(n5685), .Y(n7142) );
  CLKINVXL U9129 ( .A(w_in7[3]), .Y(n5578) );
  OAI22X1 U9130 ( .A0(n5397), .A1(n5579), .B0(n5441), .B1(n5689), .Y(n7141) );
  CLKINVXL U9131 ( .A(w_in7[4]), .Y(n5579) );
  OAI22X1 U9132 ( .A0(n5397), .A1(n5580), .B0(n5441), .B1(n5693), .Y(n7140) );
  CLKINVXL U9133 ( .A(w_in7[5]), .Y(n5580) );
  OAI22X1 U9134 ( .A0(n5396), .A1(n5581), .B0(n5441), .B1(n5697), .Y(n7139) );
  CLKINVXL U9135 ( .A(w_in7[6]), .Y(n5581) );
  OAI22X1 U9136 ( .A0(n5397), .A1(n5582), .B0(n5441), .B1(n5701), .Y(n7138) );
  CLKINVXL U9137 ( .A(w_in7[7]), .Y(n5582) );
  OAI22X1 U9138 ( .A0(n5396), .A1(n5583), .B0(n5441), .B1(n5705), .Y(n7137) );
  CLKINVXL U9139 ( .A(w_in7[8]), .Y(n5583) );
  OAI22X1 U9140 ( .A0(n5396), .A1(n5584), .B0(n5441), .B1(n5709), .Y(n7136) );
  CLKINVXL U9141 ( .A(w_in7[9]), .Y(n5584) );
  AND4X2 U9142 ( .A(n4951), .B(n4899), .C(reg_length011[0]), .D(n2484), .Y(
        n2404) );
  NOR3X1 U9143 ( .A(reg_length011[3]), .B(reg_length011[5]), .C(
        reg_length011[4]), .Y(n2484) );
  INVX2 U9144 ( .A(reg_length2[3]), .Y(n7627) );
  NOR4X1 U9145 ( .A(reg_length7[5]), .B(reg_length7[4]), .C(reg_length7[3]), 
        .D(reg_length7[2]), .Y(n2513) );
  NOR3X1 U9146 ( .A(reg_length9[3]), .B(reg_length9[5]), .C(reg_length9[4]), 
        .Y(n801) );
  INVX2 U9147 ( .A(reg_length14[4]), .Y(n7540) );
  INVX2 U9148 ( .A(reg_length8[1]), .Y(n7591) );
  INVX2 U9149 ( .A(reg_length14[3]), .Y(n7539) );
  INVX2 U9150 ( .A(reg_length14[5]), .Y(n7541) );
  INVX2 U9151 ( .A(reg_length11[2]), .Y(n7564) );
  INVX2 U9152 ( .A(reg_length11[1]), .Y(n7563) );
  NAND4X1 U9153 ( .A(n4953), .B(n4900), .C(reg_length014[0]), .D(n2523), .Y(
        n2397) );
  NOR3X1 U9154 ( .A(reg_length014[3]), .B(reg_length014[5]), .C(
        reg_length014[4]), .Y(n2523) );
  NAND2X1 U9155 ( .A(count7[0]), .B(n7273), .Y(n1706) );
  OAI2BB1X1 U9156 ( .A0N(count7[0]), .A1N(n1712), .B0(n1706), .Y(n1709) );
  OAI32X1 U9157 ( .A0(n7386), .A1(count7[2]), .A2(n1706), .B0(n1707), .B1(
        n7387), .Y(n3568) );
  AND2X1 U9158 ( .A(n1709), .B(count7[1]), .Y(n1707) );
  INVX2 U9159 ( .A(reg_length04[2]), .Y(n7409) );
  INVX2 U9160 ( .A(N5118), .Y(n5567) );
  NAND4X1 U9161 ( .A(n7573), .B(n7574), .C(N7835), .D(n808), .Y(n804) );
  NOR3X1 U9162 ( .A(reg_length10[3]), .B(reg_length10[5]), .C(reg_length10[4]), 
        .Y(n808) );
  INVX2 U9163 ( .A(reg_length04[1]), .Y(n7408) );
  OAI22X1 U9164 ( .A0(n5396), .A1(n5600), .B0(n5440), .B1(n5773), .Y(n7150) );
  OAI22X1 U9165 ( .A0(n5398), .A1(n5628), .B0(n5437), .B1(n5758), .Y(n3109) );
  OAI22X1 U9166 ( .A0(n5398), .A1(n5630), .B0(n5437), .B1(n5766), .Y(n3107) );
  INVX2 U9167 ( .A(reg_length8[5]), .Y(n7595) );
  INVX2 U9168 ( .A(reg_length9[1]), .Y(n7582) );
  INVX2 U9169 ( .A(reg_length8[4]), .Y(n7594) );
  INVX2 U9170 ( .A(y_out_sum7[36]), .Y(n6887) );
  INVX2 U9171 ( .A(reg_length9[2]), .Y(n7583) );
  MX2XL U9172 ( .A(Q12[10]), .B(x_in1[10]), .S0(n5409), .Y(n2877) );
  MX2XL U9173 ( .A(Q12[11]), .B(x_in1[11]), .S0(n5409), .Y(n2878) );
  MX2XL U9174 ( .A(Q12[12]), .B(x_in1[12]), .S0(n5408), .Y(n2879) );
  MX2XL U9175 ( .A(Q12[13]), .B(x_in1[13]), .S0(n5408), .Y(n2880) );
  MX2XL U9176 ( .A(Q12[14]), .B(x_in1[14]), .S0(n5408), .Y(n2881) );
  MX2XL U9177 ( .A(Q12[15]), .B(x_in1[15]), .S0(n5407), .Y(n2882) );
  MX2XL U9178 ( .A(Q12[1]), .B(x_in1[1]), .S0(n5410), .Y(n2883) );
  MX2XL U9179 ( .A(Q12[3]), .B(x_in1[3]), .S0(n5411), .Y(n2885) );
  MX2XL U9180 ( .A(Q12[4]), .B(x_in1[4]), .S0(n5411), .Y(n2886) );
  MX2XL U9181 ( .A(Q12[5]), .B(x_in1[5]), .S0(n5411), .Y(n2887) );
  MX2XL U9182 ( .A(Q12[6]), .B(x_in1[6]), .S0(n5410), .Y(n2888) );
  MX2XL U9183 ( .A(Q12[7]), .B(x_in1[7]), .S0(n5410), .Y(n2889) );
  MX2XL U9184 ( .A(Q12[8]), .B(x_in1[8]), .S0(n5407), .Y(n2890) );
  MX2XL U9185 ( .A(Q12[9]), .B(x_in1[9]), .S0(n5409), .Y(n2891) );
  MX2XL U9186 ( .A(Q12[2]), .B(x_in1[2]), .S0(n5412), .Y(n2884) );
  MX2XL U9187 ( .A(Q02[9]), .B(x_in0[9]), .S0(n5409), .Y(n2875) );
  MX2XL U9188 ( .A(Q02[10]), .B(x_in0[10]), .S0(n5410), .Y(n2861) );
  MX2XL U9189 ( .A(Q02[11]), .B(x_in0[11]), .S0(n5409), .Y(n2862) );
  MX2XL U9190 ( .A(Q02[12]), .B(x_in0[12]), .S0(n5408), .Y(n2863) );
  MX2XL U9191 ( .A(Q02[1]), .B(x_in0[1]), .S0(n5407), .Y(n2867) );
  MX2XL U9192 ( .A(Q02[2]), .B(x_in0[2]), .S0(n5406), .Y(n2868) );
  MX2XL U9193 ( .A(Q02[3]), .B(x_in0[3]), .S0(n5406), .Y(n2869) );
  MX2XL U9194 ( .A(Q02[4]), .B(x_in0[4]), .S0(n5406), .Y(n2870) );
  MX2XL U9195 ( .A(Q02[5]), .B(x_in0[5]), .S0(n5405), .Y(n2871) );
  MX2XL U9196 ( .A(Q02[6]), .B(x_in0[6]), .S0(n5405), .Y(n2872) );
  MX2XL U9197 ( .A(Q02[7]), .B(x_in0[7]), .S0(n5405), .Y(n2873) );
  MX2XL U9198 ( .A(Q02[8]), .B(x_in0[8]), .S0(n5407), .Y(n2874) );
  MX2XL U9199 ( .A(Q02[0]), .B(x_in0[0]), .S0(n5410), .Y(n2860) );
  MX2XL U9200 ( .A(Q12[0]), .B(x_in1[0]), .S0(n5412), .Y(n2876) );
  NOR4X1 U9201 ( .A(reg_length4[5]), .B(reg_length4[4]), .C(reg_length4[3]), 
        .D(reg_length4[2]), .Y(n2490) );
  MX2XL U9202 ( .A(Q02[13]), .B(x_in0[13]), .S0(n5407), .Y(n2864) );
  MX2XL U9203 ( .A(Q02[14]), .B(x_in0[14]), .S0(n5406), .Y(n2865) );
  INVX2 U9204 ( .A(y_out_sum7[37]), .Y(n6889) );
  NOR2X1 U9205 ( .A(N8480), .B(n7026), .Y(n2389) );
  INVX2 U9206 ( .A(n6790), .Y(n7026) );
  INVX2 U9207 ( .A(y_out_sum13[36]), .Y(n6839) );
  INVX2 U9208 ( .A(reg_length8[3]), .Y(n7593) );
  INVX2 U9209 ( .A(store_matrix7[0]), .Y(n5673) );
  INVX2 U9210 ( .A(store_matrix7[10]), .Y(n5713) );
  INVX2 U9211 ( .A(store_matrix7[11]), .Y(n5717) );
  INVX2 U9212 ( .A(store_matrix6[9]), .Y(n5773) );
  INVX2 U9213 ( .A(store_matrix7[12]), .Y(n5721) );
  INVX2 U9214 ( .A(store_matrix7[13]), .Y(n5725) );
  INVX2 U9215 ( .A(store_matrix7[14]), .Y(n5729) );
  INVX2 U9216 ( .A(store_matrix7[15]), .Y(n5733) );
  INVX2 U9217 ( .A(store_matrix6[0]), .Y(n5737) );
  INVX2 U9218 ( .A(store_matrix6[1]), .Y(n5741) );
  INVX2 U9219 ( .A(store_matrix6[2]), .Y(n5745) );
  INVX2 U9220 ( .A(store_matrix6[3]), .Y(n5749) );
  INVX2 U9221 ( .A(store_matrix6[4]), .Y(n5753) );
  INVX2 U9222 ( .A(store_matrix6[5]), .Y(n5757) );
  INVX2 U9223 ( .A(store_matrix6[6]), .Y(n5761) );
  INVX2 U9224 ( .A(store_matrix6[7]), .Y(n5765) );
  INVX2 U9225 ( .A(store_matrix6[8]), .Y(n5769) );
  INVX2 U9226 ( .A(store_matrix6[10]), .Y(n5777) );
  INVX2 U9227 ( .A(store_matrix6[11]), .Y(n5781) );
  INVX2 U9228 ( .A(store_matrix6[12]), .Y(n5785) );
  INVX2 U9229 ( .A(store_matrix6[13]), .Y(n5789) );
  INVX2 U9230 ( .A(store_matrix7[2]), .Y(n5681) );
  INVX2 U9231 ( .A(store_matrix6[14]), .Y(n5793) );
  INVX2 U9232 ( .A(store_matrix6[15]), .Y(n5797) );
  INVX2 U9233 ( .A(store_matrix7[3]), .Y(n5685) );
  INVX2 U9234 ( .A(store_matrix7[4]), .Y(n5689) );
  INVX2 U9235 ( .A(store_matrix7[5]), .Y(n5693) );
  INVX2 U9236 ( .A(store_matrix7[6]), .Y(n5697) );
  INVX2 U9237 ( .A(store_matrix7[7]), .Y(n5701) );
  INVX2 U9238 ( .A(store_matrix7[8]), .Y(n5705) );
  INVX2 U9239 ( .A(store_matrix7[9]), .Y(n5709) );
  INVX2 U9240 ( .A(y_out_sum13[37]), .Y(n6841) );
  INVX2 U9241 ( .A(reg_length10[5]), .Y(n7577) );
  INVX2 U9242 ( .A(y_out_sum9[36]), .Y(n6863) );
  INVX2 U9243 ( .A(y_out_sum7[32]), .Y(n6881) );
  INVX2 U9244 ( .A(y_out_sum7[33]), .Y(n6882) );
  INVX2 U9245 ( .A(reg_length10[1]), .Y(n7573) );
  INVX2 U9246 ( .A(store_matrix4[5]), .Y(n5758) );
  INVX2 U9247 ( .A(store_matrix4[7]), .Y(n5766) );
  INVX2 U9248 ( .A(store_matrix5[0]), .Y(n5674) );
  INVX2 U9249 ( .A(store_matrix5[1]), .Y(n5678) );
  INVX2 U9250 ( .A(store_matrix5[2]), .Y(n5682) );
  INVX2 U9251 ( .A(store_matrix5[3]), .Y(n5686) );
  INVX2 U9252 ( .A(store_matrix5[4]), .Y(n5690) );
  INVX2 U9253 ( .A(store_matrix5[5]), .Y(n5694) );
  INVX2 U9254 ( .A(store_matrix5[6]), .Y(n5698) );
  INVX2 U9255 ( .A(store_matrix5[7]), .Y(n5702) );
  INVX2 U9256 ( .A(store_matrix5[8]), .Y(n5706) );
  INVX2 U9257 ( .A(store_matrix5[9]), .Y(n5710) );
  INVX2 U9258 ( .A(store_matrix5[10]), .Y(n5714) );
  INVX2 U9259 ( .A(store_matrix5[11]), .Y(n5718) );
  INVX2 U9260 ( .A(store_matrix5[12]), .Y(n5722) );
  INVX2 U9261 ( .A(store_matrix5[13]), .Y(n5726) );
  INVX2 U9262 ( .A(store_matrix5[14]), .Y(n5730) );
  INVX2 U9263 ( .A(store_matrix5[15]), .Y(n5734) );
  INVX2 U9264 ( .A(store_matrix4[0]), .Y(n5738) );
  INVX2 U9265 ( .A(store_matrix4[1]), .Y(n5742) );
  INVX2 U9266 ( .A(store_matrix4[2]), .Y(n5746) );
  INVX2 U9267 ( .A(store_matrix4[3]), .Y(n5750) );
  INVX2 U9268 ( .A(store_matrix4[4]), .Y(n5754) );
  INVX2 U9269 ( .A(store_matrix4[6]), .Y(n5762) );
  INVX2 U9270 ( .A(store_matrix4[8]), .Y(n5770) );
  INVX2 U9271 ( .A(store_matrix4[9]), .Y(n5774) );
  INVX2 U9272 ( .A(store_matrix4[10]), .Y(n5778) );
  INVX2 U9273 ( .A(store_matrix4[11]), .Y(n5782) );
  INVX2 U9274 ( .A(store_matrix4[12]), .Y(n5786) );
  INVX2 U9275 ( .A(store_matrix4[13]), .Y(n5790) );
  INVX2 U9276 ( .A(store_matrix4[14]), .Y(n5794) );
  INVX2 U9277 ( .A(store_matrix4[15]), .Y(n5798) );
  INVX2 U9278 ( .A(y_out_sum9[37]), .Y(n6865) );
  INVX2 U9279 ( .A(store_matrix7[1]), .Y(n5677) );
  INVX2 U9280 ( .A(reg_length01[2]), .Y(n7437) );
  INVX2 U9281 ( .A(reg_length10[3]), .Y(n7575) );
  NOR4X1 U9282 ( .A(reg_length8[5]), .B(reg_length8[4]), .C(reg_length8[3]), 
        .D(reg_length8[2]), .Y(n2488) );
  INVX2 U9283 ( .A(y_out_sum13[32]), .Y(n6833) );
  INVX2 U9284 ( .A(y_out_sum12[36]), .Y(n6815) );
  INVX2 U9285 ( .A(reg_length9[4]), .Y(n7585) );
  INVX2 U9286 ( .A(reg_length9[5]), .Y(n7586) );
  INVX2 U9287 ( .A(reg_length1[2]), .Y(n7631) );
  NOR4X1 U9288 ( .A(reg_length12[5]), .B(reg_length12[4]), .C(reg_length12[3]), 
        .D(reg_length12[2]), .Y(n2475) );
  INVX2 U9289 ( .A(reg_length10[4]), .Y(n7576) );
  INVX2 U9290 ( .A(reg_length05[2]), .Y(n7401) );
  INVX2 U9291 ( .A(y_out_sum12[37]), .Y(n6817) );
  INVX2 U9292 ( .A(reg_length01[1]), .Y(n7436) );
  INVX2 U9293 ( .A(y_out_sum13[33]), .Y(n6834) );
  INVX2 U9294 ( .A(y_out_sum9[32]), .Y(n6857) );
  INVX2 U9295 ( .A(reg_length13[2]), .Y(n7546) );
  NOR4X1 U9296 ( .A(reg_length13[5]), .B(reg_length13[4]), .C(reg_length13[3]), 
        .D(reg_length13[2]), .Y(n2511) );
  INVX2 U9297 ( .A(reg_length02[2]), .Y(n7429) );
  INVX2 U9298 ( .A(y_out_sum9[33]), .Y(n6858) );
  INVX2 U9299 ( .A(reg_length5[4]), .Y(n7612) );
  INVX2 U9300 ( .A(reg_length5[5]), .Y(n7613) );
  INVX2 U9301 ( .A(reg_length9[3]), .Y(n7584) );
  INVX2 U9302 ( .A(reg_length1[1]), .Y(n7630) );
  INVX2 U9303 ( .A(reg_length05[1]), .Y(n7400) );
  INVX2 U9304 ( .A(reg_length03[2]), .Y(n7417) );
  INVX2 U9305 ( .A(reg_length2[4]), .Y(n7628) );
  INVX2 U9306 ( .A(reg_length2[5]), .Y(n7629) );
  INVX2 U9307 ( .A(reg_length7[2]), .Y(n7601) );
  INVX2 U9308 ( .A(reg_length02[1]), .Y(n7428) );
  INVX2 U9309 ( .A(y_out_sum12[32]), .Y(n6809) );
  INVX2 U9310 ( .A(reg_length10[2]), .Y(n7574) );
  NAND2X1 U9311 ( .A(count13[0]), .B(n7289), .Y(n1395) );
  OAI32X1 U9312 ( .A0(n7517), .A1(count13[2]), .A2(n1395), .B0(n1396), .B1(
        n7519), .Y(n3238) );
  INVX2 U9313 ( .A(count13[2]), .Y(n7519) );
  AND2X1 U9314 ( .A(n1398), .B(count13[1]), .Y(n1396) );
  INVX2 U9315 ( .A(y_out_sum12[33]), .Y(n6810) );
  INVX2 U9316 ( .A(reg_length5[3]), .Y(n7611) );
  INVX2 U9317 ( .A(reg_length03[1]), .Y(n7416) );
  INVX2 U9318 ( .A(reg_length7[1]), .Y(n7600) );
  NOR4X1 U9319 ( .A(reg_length11[5]), .B(reg_length11[4]), .C(reg_length11[3]), 
        .D(reg_length11[2]), .Y(n2473) );
  INVX2 U9320 ( .A(reg_length12[5]), .Y(n7558) );
  INVX2 U9321 ( .A(reg_length12[3]), .Y(n7556) );
  NAND2X1 U9322 ( .A(count8[0]), .B(n7278), .Y(n1654) );
  OAI2BB1X1 U9323 ( .A0N(count8[0]), .A1N(n1660), .B0(n1654), .Y(n1657) );
  OAI32X1 U9324 ( .A0(n7511), .A1(count8[2]), .A2(n1654), .B0(n1655), .B1(
        n7512), .Y(n3513) );
  AND2X1 U9325 ( .A(n1657), .B(count8[1]), .Y(n1655) );
  NAND2X1 U9326 ( .A(count14[0]), .B(n1350), .Y(n1342) );
  OAI32X1 U9327 ( .A0(n7504), .A1(count14[2]), .A2(n1342), .B0(n1343), .B1(
        n7505), .Y(n3183) );
  INVX2 U9328 ( .A(count14[2]), .Y(n7505) );
  AND2X1 U9329 ( .A(n1345), .B(count14[1]), .Y(n1343) );
  INVX2 U9330 ( .A(reg_length0[1]), .Y(n6788) );
  NAND2X1 U9331 ( .A(count12[0]), .B(n7280), .Y(n1449) );
  OAI2BB1X1 U9332 ( .A0N(count12[0]), .A1N(n1455), .B0(n1449), .Y(n1452) );
  OAI32X1 U9333 ( .A0(n7508), .A1(count12[2]), .A2(n1449), .B0(n1450), .B1(
        n7509), .Y(n3293) );
  AND2X1 U9334 ( .A(n1452), .B(count12[1]), .Y(n1450) );
  NAND2X1 U9335 ( .A(count10[0]), .B(n1555), .Y(n1550) );
  OAI2BB1X1 U9336 ( .A0N(count10[0]), .A1N(n1556), .B0(n1550), .Y(n1553) );
  OAI32X1 U9337 ( .A0(n7495), .A1(count10[2]), .A2(n1550), .B0(n1551), .B1(
        n7496), .Y(n3403) );
  AND2X1 U9338 ( .A(n1553), .B(count10[1]), .Y(n1551) );
  NAND2X1 U9339 ( .A(count9[0]), .B(n7288), .Y(n1601) );
  OAI2BB1X1 U9340 ( .A0N(count9[0]), .A1N(n1607), .B0(n1601), .Y(n1604) );
  OAI32X1 U9341 ( .A0(n7521), .A1(count9[2]), .A2(n1601), .B0(n1602), .B1(
        n7522), .Y(n3458) );
  AND2X1 U9342 ( .A(n1604), .B(count9[1]), .Y(n1602) );
  NAND2X1 U9343 ( .A(count6[0]), .B(n7263), .Y(n1766) );
  OAI2BB1X1 U9344 ( .A0N(count6[0]), .A1N(n1772), .B0(n1766), .Y(n1769) );
  OAI32X1 U9345 ( .A0(n7498), .A1(count6[2]), .A2(n1766), .B0(n1767), .B1(
        n7499), .Y(n3623) );
  AND2X1 U9346 ( .A(n1769), .B(count6[1]), .Y(n1767) );
  NAND2X1 U9347 ( .A(count3[0]), .B(n7274), .Y(n2015) );
  OAI2BB1X1 U9348 ( .A0N(count3[0]), .A1N(n2021), .B0(n2015), .Y(n2018) );
  OAI32X1 U9349 ( .A0(n7419), .A1(count3[2]), .A2(n2015), .B0(n2016), .B1(
        n7420), .Y(n3788) );
  AND2X1 U9350 ( .A(n2018), .B(count3[1]), .Y(n2016) );
  INVX2 U9351 ( .A(length9[2]), .Y(n7355) );
  NOR4X1 U9352 ( .A(reg_length6[5]), .B(reg_length6[4]), .C(reg_length6[3]), 
        .D(reg_length6[2]), .Y(n2509) );
  OAI32X1 U9353 ( .A0(n7385), .A1(n7273), .A2(n1712), .B0(count7[0]), .B1(
        n1713), .Y(n3569) );
  OR2X1 U9354 ( .A(n7298), .B(current_state[0]), .Y(n1314) );
  INVX2 U9355 ( .A(current_state[1]), .Y(n7298) );
  NAND2X1 U9356 ( .A(count11[0]), .B(n7271), .Y(n1501) );
  OAI2BB1X1 U9357 ( .A0N(count11[0]), .A1N(n1507), .B0(n1501), .Y(n1504) );
  OAI32X1 U9358 ( .A0(n7377), .A1(count11[2]), .A2(n1501), .B0(n1502), .B1(
        n7378), .Y(n3348) );
  AND2X1 U9359 ( .A(n1504), .B(count11[1]), .Y(n1502) );
  INVX2 U9360 ( .A(length7[2]), .Y(n7382) );
  INVX2 U9361 ( .A(length11[2]), .Y(n7373) );
  INVX2 U9362 ( .A(length12[2]), .Y(n7367) );
  INVX2 U9363 ( .A(length8[2]), .Y(n7361) );
  INVX2 U9364 ( .A(length13[2]), .Y(n7343) );
  INVX2 U9365 ( .A(length14[2]), .Y(n7337) );
  INVX2 U9366 ( .A(length10[2]), .Y(n7349) );
  OAI22X1 U9367 ( .A0(n7386), .A1(n1709), .B0(count7[1]), .B1(n1706), .Y(n3570) );
  NAND2X1 U9368 ( .A(count1[0]), .B(n7284), .Y(n2267) );
  OAI32X1 U9369 ( .A0(n7527), .A1(count1[2]), .A2(n2267), .B0(n2268), .B1(
        n7528), .Y(n3979) );
  INVX2 U9370 ( .A(count1[2]), .Y(n7528) );
  AND2X1 U9371 ( .A(n2270), .B(count1[1]), .Y(n2268) );
  NOR4X1 U9372 ( .A(n2411), .B(reg_length14[3]), .C(reg_length14[5]), .D(
        reg_length14[4]), .Y(n2410) );
  NAND2X1 U9373 ( .A(n7537), .B(n7538), .Y(n2411) );
  INVX2 U9374 ( .A(reg_length14[2]), .Y(n7538) );
  NAND2X1 U9375 ( .A(count4[0]), .B(n7276), .Y(n1933) );
  OAI2BB1X1 U9376 ( .A0N(count4[0]), .A1N(n1939), .B0(n1933), .Y(n1936) );
  OAI32X1 U9377 ( .A0(n7514), .A1(count4[2]), .A2(n1933), .B0(n1934), .B1(
        n7515), .Y(n3733) );
  AND2X1 U9378 ( .A(n1936), .B(count4[1]), .Y(n1934) );
  INVX2 U9379 ( .A(n1346), .Y(n7268) );
  AOI32X1 U9380 ( .A0(count14[0]), .A1(n7269), .A2(n1348), .B0(n7503), .B1(
        n1350), .Y(n1346) );
  INVX2 U9381 ( .A(reg_length14[1]), .Y(n7537) );
  NOR3X1 U9382 ( .A(n2263), .B(n2264), .C(n2265), .Y(n3978) );
  OAI22X1 U9383 ( .A0(n111), .A1(n171), .B0(out_valid), .B1(n5006), .Y(n2263)
         );
  INVX2 U9384 ( .A(n6791), .Y(n2264) );
  NAND4X1 U9385 ( .A(n7300), .B(n7307), .C(n114), .D(n115), .Y(n93) );
  NOR4X1 U9386 ( .A(count[15]), .B(count[13]), .C(n5378), .D(n116), .Y(n115)
         );
  AOI22X1 U9387 ( .A0(n5377), .A1(n118), .B0(count[14]), .B1(n119), .Y(n114)
         );
  AOI211X1 U9388 ( .A0(N5118), .A1(n117), .B0(count[14]), .C0(n5377), .Y(n116)
         );
  NAND2X1 U9389 ( .A(count13[2]), .B(count13[1]), .Y(n1403) );
  NAND2X1 U9390 ( .A(count5[0]), .B(n1856), .Y(n1851) );
  OAI2BB1X1 U9391 ( .A0N(count5[0]), .A1N(n1857), .B0(n1851), .Y(n1854) );
  OAI32X1 U9392 ( .A0(n7524), .A1(count5[2]), .A2(n1851), .B0(n1852), .B1(
        n7525), .Y(n3678) );
  AND2X1 U9393 ( .A(n1854), .B(count5[1]), .Y(n1852) );
  INVX2 U9394 ( .A(count12[1]), .Y(n7508) );
  INVX2 U9395 ( .A(length1[2]), .Y(n7433) );
  INVX2 U9396 ( .A(length3[2]), .Y(n7413) );
  INVX2 U9397 ( .A(length4[2]), .Y(n7405) );
  INVX2 U9398 ( .A(length5[2]), .Y(n7397) );
  INVX2 U9399 ( .A(length6[2]), .Y(n7391) );
  INVX2 U9400 ( .A(length2[2]), .Y(n7424) );
  INVX2 U9401 ( .A(count4[1]), .Y(n7514) );
  OAI32X1 U9402 ( .A0(n7418), .A1(n7274), .A2(n2021), .B0(count3[0]), .B1(
        n2022), .Y(n3789) );
  INVX2 U9403 ( .A(count6[1]), .Y(n7498) );
  INVX2 U9404 ( .A(reg_length12[4]), .Y(n7557) );
  INVX2 U9405 ( .A(count2[1]), .Y(n7501) );
  NAND2X1 U9406 ( .A(count14[2]), .B(count14[1]), .Y(n1348) );
  INVX2 U9407 ( .A(count8[1]), .Y(n7511) );
  INVX2 U9408 ( .A(count10[1]), .Y(n7495) );
  INVX2 U9409 ( .A(count13[0]), .Y(n7516) );
  INVX2 U9410 ( .A(count4[0]), .Y(n7513) );
  INVX2 U9411 ( .A(count10[0]), .Y(n7494) );
  NAND2X1 U9412 ( .A(count2[0]), .B(n2099), .Y(n2094) );
  OAI2BB1X1 U9413 ( .A0N(count2[0]), .A1N(n2100), .B0(n2094), .Y(n2097) );
  OAI32X1 U9414 ( .A0(n7501), .A1(count2[2]), .A2(n2094), .B0(n2095), .B1(
        n7502), .Y(n3843) );
  AND2X1 U9415 ( .A(n2097), .B(count2[1]), .Y(n2095) );
  INVX2 U9416 ( .A(count6[0]), .Y(n7497) );
  OAI32X1 U9417 ( .A0(n7516), .A1(n7289), .A2(n7518), .B0(count13[0]), .B1(
        n1402), .Y(n3239) );
  INVX2 U9418 ( .A(count3[1]), .Y(n7419) );
  OAI22X1 U9419 ( .A0(n7517), .A1(n1398), .B0(count13[1]), .B1(n1395), .Y(
        n3240) );
  INVX2 U9420 ( .A(n2271), .Y(n7283) );
  AOI32X1 U9421 ( .A0(count1[0]), .A1(n2272), .A2(n2273), .B0(n7526), .B1(
        n7284), .Y(n2271) );
  INVX2 U9422 ( .A(count8[0]), .Y(n7510) );
  INVX2 U9423 ( .A(count5[1]), .Y(n7524) );
  INVX2 U9424 ( .A(count2[0]), .Y(n7500) );
  INVX2 U9425 ( .A(count7[1]), .Y(n7386) );
  INVX2 U9426 ( .A(count9[1]), .Y(n7521) );
  INVX2 U9427 ( .A(count12[2]), .Y(n7509) );
  INVX2 U9428 ( .A(count4[2]), .Y(n7515) );
  INVX2 U9429 ( .A(count3[0]), .Y(n7418) );
  INVX2 U9430 ( .A(count11[1]), .Y(n7377) );
  INVX2 U9431 ( .A(count9[0]), .Y(n7520) );
  OAI32X1 U9432 ( .A0(n7510), .A1(n7278), .A2(n1660), .B0(count8[0]), .B1(
        n1661), .Y(n3514) );
  INVX2 U9433 ( .A(count11[0]), .Y(n7376) );
  INVX2 U9434 ( .A(length9[3]), .Y(n7352) );
  INVX2 U9435 ( .A(count10[2]), .Y(n7496) );
  INVX2 U9436 ( .A(count6[2]), .Y(n7499) );
  INVX2 U9437 ( .A(count5[0]), .Y(n7523) );
  INVX2 U9438 ( .A(count2[2]), .Y(n7502) );
  INVX2 U9439 ( .A(length7[3]), .Y(n7379) );
  INVX2 U9440 ( .A(length10[3]), .Y(n7346) );
  INVX2 U9441 ( .A(length11[3]), .Y(n7370) );
  INVX2 U9442 ( .A(length12[3]), .Y(n7364) );
  INVX2 U9443 ( .A(length8[3]), .Y(n7358) );
  INVX2 U9444 ( .A(length13[3]), .Y(n7340) );
  INVX2 U9445 ( .A(length14[3]), .Y(n7334) );
  OAI32X1 U9446 ( .A0(n7494), .A1(n1555), .A2(n1556), .B0(count10[0]), .B1(
        n7266), .Y(n3404) );
  INVX2 U9447 ( .A(n1555), .Y(n7266) );
  OAI22X1 U9448 ( .A0(n7511), .A1(n1657), .B0(count8[1]), .B1(n1654), .Y(n3515) );
  OAI22X1 U9449 ( .A0(n7504), .A1(n1345), .B0(count14[1]), .B1(n1342), .Y(
        n3185) );
  INVX2 U9450 ( .A(count8[2]), .Y(n7512) );
  BUFX2 U9451 ( .A(N5119), .Y(n5378) );
  INVX2 U9452 ( .A(count7[0]), .Y(n7385) );
  OAI32X1 U9453 ( .A0(n7506), .A1(n7280), .A2(n1455), .B0(count12[0]), .B1(
        n1456), .Y(n3294) );
  INVX2 U9454 ( .A(count12[0]), .Y(n7506) );
  OAI32X1 U9455 ( .A0(n7520), .A1(n7288), .A2(n1607), .B0(count9[0]), .B1(
        n1608), .Y(n3459) );
  OAI32X1 U9456 ( .A0(n7497), .A1(n7263), .A2(n1772), .B0(count6[0]), .B1(
        n1773), .Y(n3624) );
  OAI22X1 U9457 ( .A0(n7508), .A1(n1452), .B0(count12[1]), .B1(n1449), .Y(
        n3295) );
  INVX2 U9458 ( .A(count3[2]), .Y(n7420) );
  OAI22X1 U9459 ( .A0(n7495), .A1(n1553), .B0(count10[1]), .B1(n1550), .Y(
        n3405) );
  OAI22X1 U9460 ( .A0(n7521), .A1(n1604), .B0(count9[1]), .B1(n1601), .Y(n3460) );
  OAI22X1 U9461 ( .A0(n7498), .A1(n1769), .B0(count6[1]), .B1(n1766), .Y(n3625) );
  OAI32X1 U9462 ( .A0(n7513), .A1(n7276), .A2(n1939), .B0(count4[0]), .B1(
        n1940), .Y(n3734) );
  OAI32X1 U9463 ( .A0(n7376), .A1(n7271), .A2(n1507), .B0(count11[0]), .B1(
        n1508), .Y(n3349) );
  INVX2 U9464 ( .A(count5[2]), .Y(n7525) );
  INVX2 U9465 ( .A(count9[2]), .Y(n7522) );
  INVX2 U9466 ( .A(count11[2]), .Y(n7378) );
  OAI22X1 U9467 ( .A0(n7377), .A1(n1504), .B0(count11[1]), .B1(n1501), .Y(
        n3350) );
  INVX2 U9468 ( .A(count7[2]), .Y(n7387) );
  OAI32X1 U9469 ( .A0(n7500), .A1(n2099), .A2(n2100), .B0(count2[0]), .B1(
        n7262), .Y(n3844) );
  INVX2 U9470 ( .A(n2099), .Y(n7262) );
  OAI22X1 U9471 ( .A0(n7419), .A1(n2018), .B0(count3[1]), .B1(n2015), .Y(n3790) );
  OAI22X1 U9472 ( .A0(n7514), .A1(n1936), .B0(count4[1]), .B1(n1933), .Y(n3735) );
  INVX2 U9473 ( .A(length5[3]), .Y(n7394) );
  INVX2 U9474 ( .A(length1[3]), .Y(n7430) );
  INVX2 U9475 ( .A(length2[3]), .Y(n7421) );
  INVX2 U9476 ( .A(length3[3]), .Y(n7410) );
  INVX2 U9477 ( .A(length4[3]), .Y(n7402) );
  INVX2 U9478 ( .A(length6[3]), .Y(n7388) );
  ADDHXL U9479 ( .A(count_state_idle[1]), .B(count_state_idle[0]), .CO(
        r889_carry[2]), .S(N4522) );
  ADDHXL U9480 ( .A(count_state_idle[3]), .B(r889_carry[3]), .CO(r889_carry[4]), .S(N4524) );
  ADDHXL U9481 ( .A(count_state_idle[2]), .B(r889_carry[2]), .CO(r889_carry[3]), .S(N4523) );
  ADDHXL U9482 ( .A(count_state_idle[4]), .B(r889_carry[4]), .CO(r889_carry[5]), .S(N4525) );
  OAI22X1 U9483 ( .A0(n7527), .A1(n2270), .B0(count1[1]), .B1(n2267), .Y(n3981) );
  OAI32X1 U9484 ( .A0(n7523), .A1(n1856), .A2(n1857), .B0(count5[0]), .B1(
        n7287), .Y(n3679) );
  INVX2 U9485 ( .A(n1856), .Y(n7287) );
  OAI22X1 U9486 ( .A0(n7524), .A1(n1854), .B0(count5[1]), .B1(n1851), .Y(n3680) );
  INVX2 U9487 ( .A(count[13]), .Y(n7313) );
  OAI22X1 U9488 ( .A0(n7501), .A1(n2097), .B0(count2[1]), .B1(n2094), .Y(n3845) );
  BUFX2 U9489 ( .A(count[12]), .Y(n5377) );
  NOR2X1 U9490 ( .A(current_state[1]), .B(current_state[0]), .Y(n102) );
  NAND2X1 U9491 ( .A(count1[2]), .B(count1[1]), .Y(n2273) );
  BUFX2 U9492 ( .A(A3[0]), .Y(n5366) );
  BUFX2 U9493 ( .A(A3[2]), .Y(n5371) );
  BUFX2 U9494 ( .A(A3[1]), .Y(n5372) );
  INVX2 U9495 ( .A(count[15]), .Y(n7315) );
  BUFX2 U9496 ( .A(A3[5]), .Y(n5368) );
  BUFX2 U9497 ( .A(A3[4]), .Y(n5369) );
  BUFX2 U9498 ( .A(A3[3]), .Y(n5370) );
  NAND2X1 U9499 ( .A(current_state[0]), .B(n7298), .Y(N11045) );
  INVX2 U9500 ( .A(count58[5]), .Y(n7478) );
  INVX2 U9501 ( .A(count58[4]), .Y(n7477) );
  INVX2 U9502 ( .A(count58[3]), .Y(n7476) );
  INVX2 U9503 ( .A(count38[5]), .Y(n7464) );
  INVX2 U9504 ( .A(count38[4]), .Y(n7463) );
  INVX2 U9505 ( .A(count38[3]), .Y(n7462) );
  INVX2 U9506 ( .A(count1[0]), .Y(n7526) );
  INVX2 U9507 ( .A(count14[0]), .Y(n7503) );
  INVX2 U9508 ( .A(count48[5]), .Y(n7471) );
  INVX2 U9509 ( .A(count48[4]), .Y(n7470) );
  INVX2 U9510 ( .A(count48[3]), .Y(n7469) );
  INVX2 U9511 ( .A(count58[6]), .Y(n7479) );
  INVX2 U9512 ( .A(count38[6]), .Y(n7465) );
  BUFX2 U9513 ( .A(A3[6]), .Y(n5367) );
  INVX2 U9514 ( .A(count48[6]), .Y(n7472) );
  INVX2 U9515 ( .A(count08[0]), .Y(n7438) );
  INVX2 U9516 ( .A(temp_i_mat_idx[1]), .Y(n7235) );
  INVX2 U9517 ( .A(temp_i_mat_idx[0]), .Y(n7234) );
  INVX2 U9518 ( .A(count18[0]), .Y(n7445) );
  INVX2 U9519 ( .A(temp_i_mat_idx[2]), .Y(n7236) );
  INVX2 U9520 ( .A(count1[1]), .Y(n7527) );
  INVX2 U9521 ( .A(count13[1]), .Y(n7517) );
  INVX2 U9522 ( .A(count14[1]), .Y(n7504) );
  INVX2 U9523 ( .A(temp_w_mat_idx[0]), .Y(n7237) );
  INVX2 U9524 ( .A(temp_w_mat_idx[2]), .Y(n7239) );
  INVX2 U9525 ( .A(temp_w_mat_idx[1]), .Y(n7238) );
  AOI2BB2X1 U9526 ( .B0(y_out_sum9[39]), .B1(n6860), .A0N(n534), .A1N(n6859), 
        .Y(n6861) );
  OAI22X1 U9527 ( .A0(y_out_sum1[35]), .A1(n5076), .B0(y_out_sum1[33]), .B1(
        N7476), .Y(n5031) );
  OAI22X1 U9528 ( .A0(y_out_sum1[34]), .A1(n5076), .B0(y_out_sum1[32]), .B1(
        N7476), .Y(n5030) );
  AOI221XL U9529 ( .A0(n5031), .A1(N7475), .B0(n5030), .B1(reg_length1[0]), 
        .C0(N7477), .Y(n5035) );
  OAI22X1 U9530 ( .A0(y_out_sum1[38]), .A1(n5076), .B0(y_out_sum1[36]), .B1(
        N7476), .Y(n5033) );
  OAI22X1 U9531 ( .A0(y_out_sum1[39]), .A1(n5076), .B0(y_out_sum1[37]), .B1(
        N7476), .Y(n5032) );
  AOI221XL U9532 ( .A0(n5033), .A1(reg_length1[0]), .B0(N7475), .B1(n5032), 
        .C0(n5075), .Y(n5034) );
  NOR2X1 U9533 ( .A(n5035), .B(n5034), .Y(n5071) );
  NAND2X1 U9534 ( .A(N7478), .B(n5076), .Y(n5059) );
  NAND2X1 U9535 ( .A(n5074), .B(n5076), .Y(n5058) );
  OAI22X1 U9536 ( .A0(y_out_sum1[25]), .A1(n5059), .B0(y_out_sum1[17]), .B1(
        n5058), .Y(n5037) );
  NAND2X1 U9537 ( .A(N7478), .B(N7476), .Y(n5061) );
  NAND2X1 U9538 ( .A(N7476), .B(n5074), .Y(n5060) );
  OAI22X1 U9539 ( .A0(y_out_sum1[27]), .A1(n5061), .B0(y_out_sum1[19]), .B1(
        n5060), .Y(n5036) );
  NOR2X1 U9540 ( .A(n5037), .B(n5036), .Y(n5041) );
  OAI22X1 U9541 ( .A0(y_out_sum1[24]), .A1(n5059), .B0(y_out_sum1[16]), .B1(
        n5058), .Y(n5039) );
  OAI22X1 U9542 ( .A0(y_out_sum1[26]), .A1(n5061), .B0(y_out_sum1[18]), .B1(
        n5060), .Y(n5038) );
  NOR2X1 U9543 ( .A(n5039), .B(n5038), .Y(n5040) );
  OAI22X1 U9544 ( .A0(reg_length1[0]), .A1(n5041), .B0(N7475), .B1(n5040), .Y(
        n5049) );
  OAI22X1 U9545 ( .A0(y_out_sum1[29]), .A1(n5059), .B0(y_out_sum1[21]), .B1(
        n5058), .Y(n5043) );
  OAI22X1 U9546 ( .A0(y_out_sum1[31]), .A1(n5061), .B0(y_out_sum1[23]), .B1(
        n5060), .Y(n5042) );
  NOR2X1 U9547 ( .A(n5043), .B(n5042), .Y(n5047) );
  OAI22X1 U9548 ( .A0(y_out_sum1[28]), .A1(n5059), .B0(y_out_sum1[20]), .B1(
        n5058), .Y(n5045) );
  OAI22X1 U9549 ( .A0(y_out_sum1[30]), .A1(n5061), .B0(y_out_sum1[22]), .B1(
        n5060), .Y(n5044) );
  NOR2X1 U9550 ( .A(n5045), .B(n5044), .Y(n5046) );
  OAI22X1 U9551 ( .A0(reg_length1[0]), .A1(n5047), .B0(N7475), .B1(n5046), .Y(
        n5048) );
  AOI221XL U9552 ( .A0(n5049), .A1(n5075), .B0(n5048), .B1(N7477), .C0(n5072), 
        .Y(n5069) );
  OAI22X1 U9553 ( .A0(y_out_sum1[13]), .A1(n5059), .B0(y_out_sum1[5]), .B1(
        n5058), .Y(n5051) );
  OAI22X1 U9554 ( .A0(y_out_sum1[15]), .A1(n5061), .B0(y_out_sum1[7]), .B1(
        n5060), .Y(n5050) );
  NOR2X1 U9555 ( .A(n5051), .B(n5050), .Y(n5055) );
  OAI22X1 U9556 ( .A0(y_out_sum1[12]), .A1(n5059), .B0(y_out_sum1[4]), .B1(
        n5058), .Y(n5053) );
  OAI22X1 U9557 ( .A0(y_out_sum1[14]), .A1(n5061), .B0(y_out_sum1[6]), .B1(
        n5060), .Y(n5052) );
  NOR2X1 U9558 ( .A(n5053), .B(n5052), .Y(n5054) );
  OAI22X1 U9559 ( .A0(reg_length1[0]), .A1(n5055), .B0(N7475), .B1(n5054), .Y(
        n5067) );
  OAI22X1 U9560 ( .A0(y_out_sum1[9]), .A1(n5059), .B0(y_out_sum1[1]), .B1(
        n5058), .Y(n5057) );
  OAI22X1 U9561 ( .A0(y_out_sum1[11]), .A1(n5061), .B0(y_out_sum1[3]), .B1(
        n5060), .Y(n5056) );
  NOR2X1 U9562 ( .A(n5057), .B(n5056), .Y(n5065) );
  OAI22X1 U9563 ( .A0(y_out_sum1[8]), .A1(n5059), .B0(y_out_sum1[0]), .B1(
        n5058), .Y(n5063) );
  OAI22X1 U9564 ( .A0(y_out_sum1[10]), .A1(n5061), .B0(y_out_sum1[2]), .B1(
        n5060), .Y(n5062) );
  NOR2X1 U9565 ( .A(n5063), .B(n5062), .Y(n5064) );
  OAI22X1 U9566 ( .A0(reg_length1[0]), .A1(n5065), .B0(N7475), .B1(n5064), .Y(
        n5066) );
  AOI221XL U9567 ( .A0(n5067), .A1(N7477), .B0(n5066), .B1(n5075), .C0(N7479), 
        .Y(n5068) );
  NOR2X1 U9568 ( .A(n5069), .B(n5068), .Y(n5070) );
  OAI22X1 U9569 ( .A0(n5071), .A1(n5073), .B0(N7480), .B1(n5070), .Y(N9661) );
  OAI22X1 U9570 ( .A0(y_out_sum2[35]), .A1(n5121), .B0(y_out_sum2[33]), .B1(
        N7522), .Y(n5078) );
  OAI22X1 U9571 ( .A0(y_out_sum2[34]), .A1(n5121), .B0(y_out_sum2[32]), .B1(
        N7522), .Y(n5077) );
  AOI221XL U9572 ( .A0(n5078), .A1(N7521), .B0(n5077), .B1(reg_length2[0]), 
        .C0(N7523), .Y(n5082) );
  OAI22X1 U9573 ( .A0(y_out_sum2[38]), .A1(n5121), .B0(y_out_sum2[36]), .B1(
        N7522), .Y(n5080) );
  OAI22X1 U9574 ( .A0(y_out_sum2[39]), .A1(n5121), .B0(y_out_sum2[37]), .B1(
        N7522), .Y(n5079) );
  AOI221XL U9575 ( .A0(n5080), .A1(reg_length2[0]), .B0(N7521), .B1(n5079), 
        .C0(n5120), .Y(n5081) );
  NAND2X1 U9576 ( .A(N7524), .B(n5121), .Y(n5106) );
  NAND2X1 U9577 ( .A(n5119), .B(n5121), .Y(n5105) );
  OAI22X1 U9578 ( .A0(y_out_sum2[25]), .A1(n5106), .B0(y_out_sum2[17]), .B1(
        n5105), .Y(n5084) );
  NAND2X1 U9579 ( .A(N7524), .B(N7522), .Y(n5108) );
  NAND2X1 U9580 ( .A(N7522), .B(n5119), .Y(n5107) );
  OAI22X1 U9581 ( .A0(y_out_sum2[27]), .A1(n5108), .B0(y_out_sum2[19]), .B1(
        n5107), .Y(n5083) );
  NOR2X1 U9582 ( .A(n5084), .B(n5083), .Y(n5088) );
  OAI22X1 U9583 ( .A0(y_out_sum2[24]), .A1(n5106), .B0(y_out_sum2[16]), .B1(
        n5105), .Y(n5086) );
  OAI22X1 U9584 ( .A0(y_out_sum2[26]), .A1(n5108), .B0(y_out_sum2[18]), .B1(
        n5107), .Y(n5085) );
  NOR2X1 U9585 ( .A(n5086), .B(n5085), .Y(n5087) );
  OAI22X1 U9586 ( .A0(reg_length2[0]), .A1(n5088), .B0(N7521), .B1(n5087), .Y(
        n5096) );
  OAI22X1 U9587 ( .A0(y_out_sum2[29]), .A1(n5106), .B0(y_out_sum2[21]), .B1(
        n5105), .Y(n5090) );
  OAI22X1 U9588 ( .A0(y_out_sum2[31]), .A1(n5108), .B0(y_out_sum2[23]), .B1(
        n5107), .Y(n5089) );
  NOR2X1 U9589 ( .A(n5090), .B(n5089), .Y(n5094) );
  OAI22X1 U9590 ( .A0(y_out_sum2[28]), .A1(n5106), .B0(y_out_sum2[20]), .B1(
        n5105), .Y(n5092) );
  OAI22X1 U9591 ( .A0(y_out_sum2[30]), .A1(n5108), .B0(y_out_sum2[22]), .B1(
        n5107), .Y(n5091) );
  NOR2X1 U9592 ( .A(n5092), .B(n5091), .Y(n5093) );
  OAI22X1 U9593 ( .A0(reg_length2[0]), .A1(n5094), .B0(N7521), .B1(n5093), .Y(
        n5095) );
  AOI221XL U9594 ( .A0(n5096), .A1(n5120), .B0(n5095), .B1(N7523), .C0(n5118), 
        .Y(n5116) );
  OAI22X1 U9595 ( .A0(y_out_sum2[13]), .A1(n5106), .B0(y_out_sum2[5]), .B1(
        n5105), .Y(n5098) );
  OAI22X1 U9596 ( .A0(y_out_sum2[15]), .A1(n5108), .B0(y_out_sum2[7]), .B1(
        n5107), .Y(n5097) );
  NOR2X1 U9597 ( .A(n5098), .B(n5097), .Y(n5102) );
  OAI22X1 U9598 ( .A0(y_out_sum2[12]), .A1(n5106), .B0(y_out_sum2[4]), .B1(
        n5105), .Y(n5100) );
  OAI22X1 U9599 ( .A0(y_out_sum2[14]), .A1(n5108), .B0(y_out_sum2[6]), .B1(
        n5107), .Y(n5099) );
  NOR2X1 U9600 ( .A(n5100), .B(n5099), .Y(n5101) );
  OAI22X1 U9601 ( .A0(reg_length2[0]), .A1(n5102), .B0(N7521), .B1(n5101), .Y(
        n5114) );
  OAI22X1 U9602 ( .A0(y_out_sum2[9]), .A1(n5106), .B0(y_out_sum2[1]), .B1(
        n5105), .Y(n5104) );
  OAI22X1 U9603 ( .A0(y_out_sum2[11]), .A1(n5108), .B0(y_out_sum2[3]), .B1(
        n5107), .Y(n5103) );
  NOR2X1 U9604 ( .A(n5104), .B(n5103), .Y(n5112) );
  OAI22X1 U9605 ( .A0(y_out_sum2[8]), .A1(n5106), .B0(y_out_sum2[0]), .B1(
        n5105), .Y(n5110) );
  OAI22X1 U9606 ( .A0(y_out_sum2[10]), .A1(n5108), .B0(y_out_sum2[2]), .B1(
        n5107), .Y(n5109) );
  NOR2X1 U9607 ( .A(n5110), .B(n5109), .Y(n5111) );
  OAI22X1 U9608 ( .A0(reg_length2[0]), .A1(n5112), .B0(N7521), .B1(n5111), .Y(
        n5113) );
  AOI221XL U9609 ( .A0(n5114), .A1(N7523), .B0(n5113), .B1(n5120), .C0(N7525), 
        .Y(n5115) );
  NOR2X1 U9610 ( .A(n5116), .B(n5115), .Y(n5117) );
  OAI22X1 U9611 ( .A0(y_out_sum3[35]), .A1(n5166), .B0(y_out_sum3[33]), .B1(
        N7566), .Y(n5123) );
  OAI22X1 U9612 ( .A0(y_out_sum3[34]), .A1(n5166), .B0(y_out_sum3[32]), .B1(
        N7566), .Y(n5122) );
  AOI221XL U9613 ( .A0(n5123), .A1(N7565), .B0(n5122), .B1(reg_length3[0]), 
        .C0(N7567), .Y(n5127) );
  OAI22X1 U9614 ( .A0(y_out_sum3[38]), .A1(n5166), .B0(y_out_sum3[36]), .B1(
        N7566), .Y(n5125) );
  OAI22X1 U9615 ( .A0(y_out_sum3[39]), .A1(n5166), .B0(y_out_sum3[37]), .B1(
        N7566), .Y(n5124) );
  AOI221XL U9616 ( .A0(n5125), .A1(reg_length3[0]), .B0(N7565), .B1(n5124), 
        .C0(n5165), .Y(n5126) );
  NAND2X1 U9617 ( .A(N7568), .B(n5166), .Y(n5151) );
  NAND2X1 U9618 ( .A(n5164), .B(n5166), .Y(n5150) );
  OAI22X1 U9619 ( .A0(y_out_sum3[25]), .A1(n5151), .B0(y_out_sum3[17]), .B1(
        n5150), .Y(n5129) );
  NAND2X1 U9620 ( .A(N7568), .B(N7566), .Y(n5153) );
  NAND2X1 U9621 ( .A(N7566), .B(n5164), .Y(n5152) );
  OAI22X1 U9622 ( .A0(y_out_sum3[27]), .A1(n5153), .B0(y_out_sum3[19]), .B1(
        n5152), .Y(n5128) );
  NOR2X1 U9623 ( .A(n5129), .B(n5128), .Y(n5133) );
  OAI22X1 U9624 ( .A0(y_out_sum3[24]), .A1(n5151), .B0(y_out_sum3[16]), .B1(
        n5150), .Y(n5131) );
  OAI22X1 U9625 ( .A0(y_out_sum3[26]), .A1(n5153), .B0(y_out_sum3[18]), .B1(
        n5152), .Y(n5130) );
  NOR2X1 U9626 ( .A(n5131), .B(n5130), .Y(n5132) );
  OAI22X1 U9627 ( .A0(reg_length3[0]), .A1(n5133), .B0(N7565), .B1(n5132), .Y(
        n5141) );
  OAI22X1 U9628 ( .A0(y_out_sum3[29]), .A1(n5151), .B0(y_out_sum3[21]), .B1(
        n5150), .Y(n5135) );
  OAI22X1 U9629 ( .A0(y_out_sum3[31]), .A1(n5153), .B0(y_out_sum3[23]), .B1(
        n5152), .Y(n5134) );
  NOR2X1 U9630 ( .A(n5135), .B(n5134), .Y(n5139) );
  OAI22X1 U9631 ( .A0(y_out_sum3[28]), .A1(n5151), .B0(y_out_sum3[20]), .B1(
        n5150), .Y(n5137) );
  OAI22X1 U9632 ( .A0(y_out_sum3[30]), .A1(n5153), .B0(y_out_sum3[22]), .B1(
        n5152), .Y(n5136) );
  NOR2X1 U9633 ( .A(n5137), .B(n5136), .Y(n5138) );
  OAI22X1 U9634 ( .A0(reg_length3[0]), .A1(n5139), .B0(N7565), .B1(n5138), .Y(
        n5140) );
  AOI221XL U9635 ( .A0(n5141), .A1(n5165), .B0(n5140), .B1(N7567), .C0(n5163), 
        .Y(n5161) );
  OAI22X1 U9636 ( .A0(y_out_sum3[13]), .A1(n5151), .B0(y_out_sum3[5]), .B1(
        n5150), .Y(n5143) );
  OAI22X1 U9637 ( .A0(y_out_sum3[15]), .A1(n5153), .B0(y_out_sum3[7]), .B1(
        n5152), .Y(n5142) );
  NOR2X1 U9638 ( .A(n5143), .B(n5142), .Y(n5147) );
  OAI22X1 U9639 ( .A0(y_out_sum3[12]), .A1(n5151), .B0(y_out_sum3[4]), .B1(
        n5150), .Y(n5145) );
  OAI22X1 U9640 ( .A0(y_out_sum3[14]), .A1(n5153), .B0(y_out_sum3[6]), .B1(
        n5152), .Y(n5144) );
  NOR2X1 U9641 ( .A(n5145), .B(n5144), .Y(n5146) );
  OAI22X1 U9642 ( .A0(reg_length3[0]), .A1(n5147), .B0(N7565), .B1(n5146), .Y(
        n5159) );
  OAI22X1 U9643 ( .A0(y_out_sum3[9]), .A1(n5151), .B0(y_out_sum3[1]), .B1(
        n5150), .Y(n5149) );
  OAI22X1 U9644 ( .A0(y_out_sum3[11]), .A1(n5153), .B0(y_out_sum3[3]), .B1(
        n5152), .Y(n5148) );
  NOR2X1 U9645 ( .A(n5149), .B(n5148), .Y(n5157) );
  OAI22X1 U9646 ( .A0(y_out_sum3[8]), .A1(n5151), .B0(y_out_sum3[0]), .B1(
        n5150), .Y(n5155) );
  OAI22X1 U9647 ( .A0(y_out_sum3[10]), .A1(n5153), .B0(y_out_sum3[2]), .B1(
        n5152), .Y(n5154) );
  NOR2X1 U9648 ( .A(n5155), .B(n5154), .Y(n5156) );
  OAI22X1 U9649 ( .A0(reg_length3[0]), .A1(n5157), .B0(N7565), .B1(n5156), .Y(
        n5158) );
  AOI221XL U9650 ( .A0(n5159), .A1(N7567), .B0(n5158), .B1(n5165), .C0(N7569), 
        .Y(n5160) );
  NOR2X1 U9651 ( .A(n5161), .B(n5160), .Y(n5162) );
  OAI22X1 U9652 ( .A0(y_out_sum4[35]), .A1(n5211), .B0(y_out_sum4[33]), .B1(
        N7607), .Y(n5168) );
  OAI22X1 U9653 ( .A0(y_out_sum4[34]), .A1(n5211), .B0(y_out_sum4[32]), .B1(
        N7607), .Y(n5167) );
  AOI221XL U9654 ( .A0(n5168), .A1(N7606), .B0(n5167), .B1(reg_length4[0]), 
        .C0(N7608), .Y(n5172) );
  OAI22X1 U9655 ( .A0(y_out_sum4[38]), .A1(n5211), .B0(y_out_sum4[36]), .B1(
        N7607), .Y(n5170) );
  OAI22X1 U9656 ( .A0(y_out_sum4[39]), .A1(n5211), .B0(y_out_sum4[37]), .B1(
        N7607), .Y(n5169) );
  AOI221XL U9657 ( .A0(n5170), .A1(reg_length4[0]), .B0(N7606), .B1(n5169), 
        .C0(n5210), .Y(n5171) );
  NAND2X1 U9658 ( .A(N7609), .B(n5211), .Y(n5196) );
  NAND2X1 U9659 ( .A(n5209), .B(n5211), .Y(n5195) );
  OAI22X1 U9660 ( .A0(y_out_sum4[25]), .A1(n5196), .B0(y_out_sum4[17]), .B1(
        n5195), .Y(n5174) );
  NAND2X1 U9661 ( .A(N7609), .B(N7607), .Y(n5198) );
  NAND2X1 U9662 ( .A(N7607), .B(n5209), .Y(n5197) );
  OAI22X1 U9663 ( .A0(y_out_sum4[27]), .A1(n5198), .B0(y_out_sum4[19]), .B1(
        n5197), .Y(n5173) );
  NOR2X1 U9664 ( .A(n5174), .B(n5173), .Y(n5178) );
  OAI22X1 U9665 ( .A0(y_out_sum4[24]), .A1(n5196), .B0(y_out_sum4[16]), .B1(
        n5195), .Y(n5176) );
  OAI22X1 U9666 ( .A0(y_out_sum4[26]), .A1(n5198), .B0(y_out_sum4[18]), .B1(
        n5197), .Y(n5175) );
  NOR2X1 U9667 ( .A(n5176), .B(n5175), .Y(n5177) );
  OAI22X1 U9668 ( .A0(reg_length4[0]), .A1(n5178), .B0(N7606), .B1(n5177), .Y(
        n5186) );
  OAI22X1 U9669 ( .A0(y_out_sum4[29]), .A1(n5196), .B0(y_out_sum4[21]), .B1(
        n5195), .Y(n5180) );
  OAI22X1 U9670 ( .A0(y_out_sum4[31]), .A1(n5198), .B0(y_out_sum4[23]), .B1(
        n5197), .Y(n5179) );
  NOR2X1 U9671 ( .A(n5180), .B(n5179), .Y(n5184) );
  OAI22X1 U9672 ( .A0(y_out_sum4[28]), .A1(n5196), .B0(y_out_sum4[20]), .B1(
        n5195), .Y(n5182) );
  OAI22X1 U9673 ( .A0(y_out_sum4[30]), .A1(n5198), .B0(y_out_sum4[22]), .B1(
        n5197), .Y(n5181) );
  NOR2X1 U9674 ( .A(n5182), .B(n5181), .Y(n5183) );
  OAI22X1 U9675 ( .A0(reg_length4[0]), .A1(n5184), .B0(N7606), .B1(n5183), .Y(
        n5185) );
  AOI221XL U9676 ( .A0(n5186), .A1(n5210), .B0(n5185), .B1(N7608), .C0(n5208), 
        .Y(n5206) );
  OAI22X1 U9677 ( .A0(y_out_sum4[13]), .A1(n5196), .B0(y_out_sum4[5]), .B1(
        n5195), .Y(n5188) );
  OAI22X1 U9678 ( .A0(y_out_sum4[15]), .A1(n5198), .B0(y_out_sum4[7]), .B1(
        n5197), .Y(n5187) );
  NOR2X1 U9679 ( .A(n5188), .B(n5187), .Y(n5192) );
  OAI22X1 U9680 ( .A0(y_out_sum4[12]), .A1(n5196), .B0(y_out_sum4[4]), .B1(
        n5195), .Y(n5190) );
  OAI22X1 U9681 ( .A0(y_out_sum4[14]), .A1(n5198), .B0(y_out_sum4[6]), .B1(
        n5197), .Y(n5189) );
  NOR2X1 U9682 ( .A(n5190), .B(n5189), .Y(n5191) );
  OAI22X1 U9683 ( .A0(reg_length4[0]), .A1(n5192), .B0(N7606), .B1(n5191), .Y(
        n5204) );
  OAI22X1 U9684 ( .A0(y_out_sum4[9]), .A1(n5196), .B0(y_out_sum4[1]), .B1(
        n5195), .Y(n5194) );
  OAI22X1 U9685 ( .A0(y_out_sum4[11]), .A1(n5198), .B0(y_out_sum4[3]), .B1(
        n5197), .Y(n5193) );
  NOR2X1 U9686 ( .A(n5194), .B(n5193), .Y(n5202) );
  OAI22X1 U9687 ( .A0(y_out_sum4[8]), .A1(n5196), .B0(y_out_sum4[0]), .B1(
        n5195), .Y(n5200) );
  OAI22X1 U9688 ( .A0(y_out_sum4[10]), .A1(n5198), .B0(y_out_sum4[2]), .B1(
        n5197), .Y(n5199) );
  NOR2X1 U9689 ( .A(n5200), .B(n5199), .Y(n5201) );
  OAI22X1 U9690 ( .A0(reg_length4[0]), .A1(n5202), .B0(N7606), .B1(n5201), .Y(
        n5203) );
  AOI221XL U9691 ( .A0(n5204), .A1(N7608), .B0(n5203), .B1(n5210), .C0(N7610), 
        .Y(n5205) );
  NOR2X1 U9692 ( .A(n5206), .B(n5205), .Y(n5207) );
  OAI22X1 U9693 ( .A0(y_out_sum5[35]), .A1(n5256), .B0(y_out_sum5[33]), .B1(
        N7648), .Y(n5213) );
  OAI22X1 U9694 ( .A0(y_out_sum5[34]), .A1(n5256), .B0(y_out_sum5[32]), .B1(
        N7648), .Y(n5212) );
  AOI221XL U9695 ( .A0(n5213), .A1(n4934), .B0(n5212), .B1(reg_length5[0]), 
        .C0(N7649), .Y(n5217) );
  OAI22X1 U9696 ( .A0(y_out_sum5[38]), .A1(n5256), .B0(y_out_sum5[36]), .B1(
        N7648), .Y(n5215) );
  OAI22X1 U9697 ( .A0(y_out_sum5[39]), .A1(n5256), .B0(y_out_sum5[37]), .B1(
        N7648), .Y(n5214) );
  AOI221XL U9698 ( .A0(n5215), .A1(reg_length5[0]), .B0(n4934), .B1(n5214), 
        .C0(n5255), .Y(n5216) );
  NAND2X1 U9699 ( .A(N7650), .B(n5256), .Y(n5241) );
  NAND2X1 U9700 ( .A(n5254), .B(n5256), .Y(n5240) );
  OAI22X1 U9701 ( .A0(y_out_sum5[25]), .A1(n5241), .B0(y_out_sum5[17]), .B1(
        n5240), .Y(n5219) );
  NAND2X1 U9702 ( .A(N7650), .B(N7648), .Y(n5243) );
  NAND2X1 U9703 ( .A(N7648), .B(n5254), .Y(n5242) );
  OAI22X1 U9704 ( .A0(y_out_sum5[27]), .A1(n5243), .B0(y_out_sum5[19]), .B1(
        n5242), .Y(n5218) );
  NOR2X1 U9705 ( .A(n5219), .B(n5218), .Y(n5223) );
  OAI22X1 U9706 ( .A0(y_out_sum5[24]), .A1(n5241), .B0(y_out_sum5[16]), .B1(
        n5240), .Y(n5221) );
  OAI22X1 U9707 ( .A0(y_out_sum5[26]), .A1(n5243), .B0(y_out_sum5[18]), .B1(
        n5242), .Y(n5220) );
  NOR2X1 U9708 ( .A(n5221), .B(n5220), .Y(n5222) );
  OAI22X1 U9709 ( .A0(reg_length5[0]), .A1(n5223), .B0(n4934), .B1(n5222), .Y(
        n5231) );
  OAI22X1 U9710 ( .A0(y_out_sum5[29]), .A1(n5241), .B0(y_out_sum5[21]), .B1(
        n5240), .Y(n5225) );
  OAI22X1 U9711 ( .A0(y_out_sum5[31]), .A1(n5243), .B0(y_out_sum5[23]), .B1(
        n5242), .Y(n5224) );
  NOR2X1 U9712 ( .A(n5225), .B(n5224), .Y(n5229) );
  OAI22X1 U9713 ( .A0(y_out_sum5[28]), .A1(n5241), .B0(y_out_sum5[20]), .B1(
        n5240), .Y(n5227) );
  OAI22X1 U9714 ( .A0(y_out_sum5[30]), .A1(n5243), .B0(y_out_sum5[22]), .B1(
        n5242), .Y(n5226) );
  NOR2X1 U9715 ( .A(n5227), .B(n5226), .Y(n5228) );
  OAI22X1 U9716 ( .A0(reg_length5[0]), .A1(n5229), .B0(n4934), .B1(n5228), .Y(
        n5230) );
  AOI221XL U9717 ( .A0(n5231), .A1(n5255), .B0(n5230), .B1(N7649), .C0(n5253), 
        .Y(n5251) );
  OAI22X1 U9718 ( .A0(y_out_sum5[13]), .A1(n5241), .B0(y_out_sum5[5]), .B1(
        n5240), .Y(n5233) );
  OAI22X1 U9719 ( .A0(y_out_sum5[15]), .A1(n5243), .B0(y_out_sum5[7]), .B1(
        n5242), .Y(n5232) );
  NOR2X1 U9720 ( .A(n5233), .B(n5232), .Y(n5237) );
  OAI22X1 U9721 ( .A0(y_out_sum5[12]), .A1(n5241), .B0(y_out_sum5[4]), .B1(
        n5240), .Y(n5235) );
  OAI22X1 U9722 ( .A0(y_out_sum5[14]), .A1(n5243), .B0(y_out_sum5[6]), .B1(
        n5242), .Y(n5234) );
  NOR2X1 U9723 ( .A(n5235), .B(n5234), .Y(n5236) );
  OAI22X1 U9724 ( .A0(reg_length5[0]), .A1(n5237), .B0(n4934), .B1(n5236), .Y(
        n5249) );
  OAI22X1 U9725 ( .A0(y_out_sum5[9]), .A1(n5241), .B0(y_out_sum5[1]), .B1(
        n5240), .Y(n5239) );
  OAI22X1 U9726 ( .A0(y_out_sum5[11]), .A1(n5243), .B0(y_out_sum5[3]), .B1(
        n5242), .Y(n5238) );
  NOR2X1 U9727 ( .A(n5239), .B(n5238), .Y(n5247) );
  OAI22X1 U9728 ( .A0(y_out_sum5[8]), .A1(n5241), .B0(y_out_sum5[0]), .B1(
        n5240), .Y(n5245) );
  OAI22X1 U9729 ( .A0(y_out_sum5[10]), .A1(n5243), .B0(y_out_sum5[2]), .B1(
        n5242), .Y(n5244) );
  NOR2X1 U9730 ( .A(n5245), .B(n5244), .Y(n5246) );
  OAI22X1 U9731 ( .A0(reg_length5[0]), .A1(n5247), .B0(n4934), .B1(n5246), .Y(
        n5248) );
  AOI221XL U9732 ( .A0(n5249), .A1(N7649), .B0(n5248), .B1(n5255), .C0(N7651), 
        .Y(n5250) );
  NOR2X1 U9733 ( .A(n5251), .B(n5250), .Y(n5252) );
  OAI22X1 U9734 ( .A0(y_out_sum6[35]), .A1(n5301), .B0(y_out_sum6[33]), .B1(
        N7689), .Y(n5258) );
  OAI22X1 U9735 ( .A0(y_out_sum6[34]), .A1(n5301), .B0(y_out_sum6[32]), .B1(
        N7689), .Y(n5257) );
  AOI221XL U9736 ( .A0(n5258), .A1(N7688), .B0(n5257), .B1(reg_length6[0]), 
        .C0(N7690), .Y(n5262) );
  OAI22X1 U9737 ( .A0(y_out_sum6[38]), .A1(n5301), .B0(y_out_sum6[36]), .B1(
        N7689), .Y(n5260) );
  OAI22X1 U9738 ( .A0(y_out_sum6[39]), .A1(n5301), .B0(y_out_sum6[37]), .B1(
        N7689), .Y(n5259) );
  AOI221XL U9739 ( .A0(n5260), .A1(reg_length6[0]), .B0(N7688), .B1(n5259), 
        .C0(n5300), .Y(n5261) );
  NAND2X1 U9740 ( .A(N7691), .B(n5301), .Y(n5286) );
  NAND2X1 U9741 ( .A(n5299), .B(n5301), .Y(n5285) );
  OAI22X1 U9742 ( .A0(y_out_sum6[25]), .A1(n5286), .B0(y_out_sum6[17]), .B1(
        n5285), .Y(n5264) );
  NAND2X1 U9743 ( .A(N7691), .B(N7689), .Y(n5288) );
  NAND2X1 U9744 ( .A(N7689), .B(n5299), .Y(n5287) );
  OAI22X1 U9745 ( .A0(y_out_sum6[27]), .A1(n5288), .B0(y_out_sum6[19]), .B1(
        n5287), .Y(n5263) );
  NOR2X1 U9746 ( .A(n5264), .B(n5263), .Y(n5268) );
  OAI22X1 U9747 ( .A0(y_out_sum6[24]), .A1(n5286), .B0(y_out_sum6[16]), .B1(
        n5285), .Y(n5266) );
  OAI22X1 U9748 ( .A0(y_out_sum6[26]), .A1(n5288), .B0(y_out_sum6[18]), .B1(
        n5287), .Y(n5265) );
  NOR2X1 U9749 ( .A(n5266), .B(n5265), .Y(n5267) );
  OAI22X1 U9750 ( .A0(reg_length6[0]), .A1(n5268), .B0(N7688), .B1(n5267), .Y(
        n5276) );
  OAI22X1 U9751 ( .A0(y_out_sum6[29]), .A1(n5286), .B0(y_out_sum6[21]), .B1(
        n5285), .Y(n5270) );
  OAI22X1 U9752 ( .A0(y_out_sum6[31]), .A1(n5288), .B0(y_out_sum6[23]), .B1(
        n5287), .Y(n5269) );
  NOR2X1 U9753 ( .A(n5270), .B(n5269), .Y(n5274) );
  OAI22X1 U9754 ( .A0(y_out_sum6[28]), .A1(n5286), .B0(y_out_sum6[20]), .B1(
        n5285), .Y(n5272) );
  OAI22X1 U9755 ( .A0(y_out_sum6[30]), .A1(n5288), .B0(y_out_sum6[22]), .B1(
        n5287), .Y(n5271) );
  NOR2X1 U9756 ( .A(n5272), .B(n5271), .Y(n5273) );
  OAI22X1 U9757 ( .A0(reg_length6[0]), .A1(n5274), .B0(N7688), .B1(n5273), .Y(
        n5275) );
  AOI221XL U9758 ( .A0(n5276), .A1(n5300), .B0(n5275), .B1(N7690), .C0(n5298), 
        .Y(n5296) );
  OAI22X1 U9759 ( .A0(y_out_sum6[13]), .A1(n5286), .B0(y_out_sum6[5]), .B1(
        n5285), .Y(n5278) );
  OAI22X1 U9760 ( .A0(y_out_sum6[15]), .A1(n5288), .B0(y_out_sum6[7]), .B1(
        n5287), .Y(n5277) );
  NOR2X1 U9761 ( .A(n5278), .B(n5277), .Y(n5282) );
  OAI22X1 U9762 ( .A0(y_out_sum6[12]), .A1(n5286), .B0(y_out_sum6[4]), .B1(
        n5285), .Y(n5280) );
  OAI22X1 U9763 ( .A0(y_out_sum6[14]), .A1(n5288), .B0(y_out_sum6[6]), .B1(
        n5287), .Y(n5279) );
  NOR2X1 U9764 ( .A(n5280), .B(n5279), .Y(n5281) );
  OAI22X1 U9765 ( .A0(reg_length6[0]), .A1(n5282), .B0(N7688), .B1(n5281), .Y(
        n5294) );
  OAI22X1 U9766 ( .A0(y_out_sum6[9]), .A1(n5286), .B0(y_out_sum6[1]), .B1(
        n5285), .Y(n5284) );
  OAI22X1 U9767 ( .A0(y_out_sum6[11]), .A1(n5288), .B0(y_out_sum6[3]), .B1(
        n5287), .Y(n5283) );
  NOR2X1 U9768 ( .A(n5284), .B(n5283), .Y(n5292) );
  OAI22X1 U9769 ( .A0(y_out_sum6[8]), .A1(n5286), .B0(y_out_sum6[0]), .B1(
        n5285), .Y(n5290) );
  OAI22X1 U9770 ( .A0(y_out_sum6[10]), .A1(n5288), .B0(y_out_sum6[2]), .B1(
        n5287), .Y(n5289) );
  NOR2X1 U9771 ( .A(n5290), .B(n5289), .Y(n5291) );
  OAI22X1 U9772 ( .A0(reg_length6[0]), .A1(n5292), .B0(N7688), .B1(n5291), .Y(
        n5293) );
  AOI221XL U9773 ( .A0(n5294), .A1(N7690), .B0(n5293), .B1(n5300), .C0(N7692), 
        .Y(n5295) );
  NOR2X1 U9774 ( .A(n5296), .B(n5295), .Y(n5297) );
  OAI22X1 U9775 ( .A0(y_out_sum0[35]), .A1(n5345), .B0(y_out_sum0[33]), .B1(
        N7430), .Y(n5303) );
  OAI22X1 U9776 ( .A0(y_out_sum0[34]), .A1(n5345), .B0(y_out_sum0[32]), .B1(
        N7430), .Y(n5302) );
  AOI221XL U9777 ( .A0(n5303), .A1(N7429), .B0(n5302), .B1(reg_length0[0]), 
        .C0(N7431), .Y(n5307) );
  OAI22X1 U9778 ( .A0(y_out_sum0[38]), .A1(n5345), .B0(y_out_sum0[36]), .B1(
        N7430), .Y(n5305) );
  OAI22X1 U9779 ( .A0(y_out_sum0[39]), .A1(n5345), .B0(y_out_sum0[37]), .B1(
        N7430), .Y(n5304) );
  AOI221XL U9780 ( .A0(n5305), .A1(reg_length0[0]), .B0(N7429), .B1(n5304), 
        .C0(n5344), .Y(n5306) );
  NOR2X1 U9781 ( .A(n5307), .B(n5306), .Y(n5343) );
  NAND2X1 U9782 ( .A(N7432), .B(n5345), .Y(n5331) );
  NAND2X1 U9783 ( .A(n5346), .B(n5345), .Y(n5330) );
  OAI22X1 U9784 ( .A0(y_out_sum0[25]), .A1(n5331), .B0(y_out_sum0[17]), .B1(
        n5330), .Y(n5309) );
  NAND2X1 U9785 ( .A(N7432), .B(N7430), .Y(n5333) );
  NAND2X1 U9786 ( .A(N7430), .B(n5346), .Y(n5332) );
  OAI22X1 U9787 ( .A0(y_out_sum0[27]), .A1(n5333), .B0(y_out_sum0[19]), .B1(
        n5332), .Y(n5308) );
  NOR2X1 U9788 ( .A(n5309), .B(n5308), .Y(n5313) );
  OAI22X1 U9789 ( .A0(y_out_sum0[24]), .A1(n5331), .B0(y_out_sum0[16]), .B1(
        n5330), .Y(n5311) );
  OAI22X1 U9790 ( .A0(y_out_sum0[26]), .A1(n5333), .B0(y_out_sum0[18]), .B1(
        n5332), .Y(n5310) );
  NOR2X1 U9791 ( .A(n5311), .B(n5310), .Y(n5312) );
  OAI22X1 U9792 ( .A0(reg_length0[0]), .A1(n5313), .B0(N7429), .B1(n5312), .Y(
        n5321) );
  OAI22X1 U9793 ( .A0(y_out_sum0[29]), .A1(n5331), .B0(y_out_sum0[21]), .B1(
        n5330), .Y(n5315) );
  OAI22X1 U9794 ( .A0(y_out_sum0[31]), .A1(n5333), .B0(y_out_sum0[23]), .B1(
        n5332), .Y(n5314) );
  NOR2X1 U9795 ( .A(n5315), .B(n5314), .Y(n5319) );
  OAI22X1 U9796 ( .A0(y_out_sum0[28]), .A1(n5331), .B0(y_out_sum0[20]), .B1(
        n5330), .Y(n5317) );
  OAI22X1 U9797 ( .A0(y_out_sum0[30]), .A1(n5333), .B0(y_out_sum0[22]), .B1(
        n5332), .Y(n5316) );
  NOR2X1 U9798 ( .A(n5317), .B(n5316), .Y(n5318) );
  OAI22X1 U9799 ( .A0(reg_length0[0]), .A1(n5319), .B0(N7429), .B1(n5318), .Y(
        n5320) );
  AOI221XL U9800 ( .A0(n5321), .A1(n5344), .B0(n5320), .B1(N7431), .C0(n6032), 
        .Y(n5341) );
  OAI22X1 U9801 ( .A0(y_out_sum0[13]), .A1(n5331), .B0(y_out_sum0[5]), .B1(
        n5330), .Y(n5323) );
  OAI22X1 U9802 ( .A0(y_out_sum0[15]), .A1(n5333), .B0(y_out_sum0[7]), .B1(
        n5332), .Y(n5322) );
  NOR2X1 U9803 ( .A(n5323), .B(n5322), .Y(n5327) );
  OAI22X1 U9804 ( .A0(y_out_sum0[12]), .A1(n5331), .B0(y_out_sum0[4]), .B1(
        n5330), .Y(n5325) );
  OAI22X1 U9805 ( .A0(y_out_sum0[14]), .A1(n5333), .B0(y_out_sum0[6]), .B1(
        n5332), .Y(n5324) );
  NOR2X1 U9806 ( .A(n5325), .B(n5324), .Y(n5326) );
  OAI22X1 U9807 ( .A0(reg_length0[0]), .A1(n5327), .B0(N7429), .B1(n5326), .Y(
        n5339) );
  OAI22X1 U9808 ( .A0(y_out_sum0[9]), .A1(n5331), .B0(y_out_sum0[1]), .B1(
        n5330), .Y(n5329) );
  OAI22X1 U9809 ( .A0(y_out_sum0[11]), .A1(n5333), .B0(y_out_sum0[3]), .B1(
        n5332), .Y(n5328) );
  NOR2X1 U9810 ( .A(n5329), .B(n5328), .Y(n5337) );
  OAI22X1 U9811 ( .A0(y_out_sum0[8]), .A1(n5331), .B0(y_out_sum0[0]), .B1(
        n5330), .Y(n5335) );
  OAI22X1 U9812 ( .A0(y_out_sum0[10]), .A1(n5333), .B0(y_out_sum0[2]), .B1(
        n5332), .Y(n5334) );
  NOR2X1 U9813 ( .A(n5335), .B(n5334), .Y(n5336) );
  OAI22X1 U9814 ( .A0(reg_length0[0]), .A1(n5337), .B0(N7429), .B1(n5336), .Y(
        n5338) );
  AOI221XL U9815 ( .A0(n5339), .A1(N7431), .B0(n5338), .B1(n5344), .C0(N7433), 
        .Y(n5340) );
  NOR2X1 U9816 ( .A(n5341), .B(n5340), .Y(n5342) );
  OAI22X1 U9817 ( .A0(n5343), .A1(n6040), .B0(N7434), .B1(n5342), .Y(N9425) );
  OAI2BB1XL U9818 ( .A0N(n5971), .A1N(n5563), .B0(n5561), .Y(n5972) );
  OAI2BB1X1 U9819 ( .A0N(n5969), .A1N(n5550), .B0(n5552), .Y(n5970) );
  CLKINVXL U9820 ( .A(sum[39]), .Y(n5558) );
  CLKINVX2 U9821 ( .A(sum[34]), .Y(n5554) );
  OAI22X1 U9822 ( .A0(n5397), .A1(n5576), .B0(n5441), .B1(n5677), .Y(n7156) );
  CLKINVXL U9823 ( .A(w_in7[1]), .Y(n5576) );
  MX2XL U9824 ( .A(Q02[15]), .B(x_in0[15]), .S0(n5405), .Y(n2866) );
  OAI2BB1XL U9825 ( .A0N(reg_length00[3]), .A1N(n6787), .B0(n6784), .Y(n3173)
         );
  MX2X2 U9826 ( .A(n7010), .B(out_value), .S0(n7009), .Y(n2859) );
  OR3X2 U9827 ( .A(reg_matrix_size[1]), .B(n7036), .C(reg_matrix_size[2]), .Y(
        n7232) );
  OR3X2 U9828 ( .A(reg_matrix_size[1]), .B(n5574), .C(reg_matrix_size[3]), .Y(
        n111) );
  OR4X2 U9829 ( .A(n5442), .B(n5899), .C(n5898), .D(n7270), .Y(n6791) );
  OR3X2 U9830 ( .A(reg_invalid2[0]), .B(n6776), .C(n6777), .Y(n2783) );
  OR3X2 U9831 ( .A(n2461), .B(n6775), .C(n96), .Y(n6790) );
  OR3X2 U9832 ( .A(n7047), .B(n96), .C(n6778), .Y(n6037) );
  OR4X2 U9833 ( .A(n5493), .B(n6009), .C(n5495), .D(n5977), .Y(n5951) );
  OR2X4 U9834 ( .A(n5549), .B(n5547), .Y(n5995) );
  OR4X2 U9835 ( .A(n5482), .B(n5485), .C(n5489), .D(n4967), .Y(n6010) );
  OR4X2 U9836 ( .A(n5531), .B(n6018), .C(n4976), .D(n6017), .Y(n6021) );
  OR3X2 U9837 ( .A(sum[23]), .B(n6028), .C(n6027), .Y(n6029) );
  OR4X2 U9838 ( .A(n7321), .B(n7022), .C(n2073), .D(n2072), .Y(n6188) );
  OR3X2 U9839 ( .A(n2697), .B(n7230), .C(n2814), .Y(n6608) );
  OR3X2 U9840 ( .A(n2461), .B(n7230), .C(n1585), .Y(n6665) );
  OR3X2 U9841 ( .A(n2805), .B(n5376), .C(n6719), .Y(n6720) );
  OR4X2 U9842 ( .A(reg_length0[2]), .B(reg_length0[3]), .C(reg_length0[5]), 
        .D(reg_length0[4]), .Y(n6789) );
  OR4X2 U9843 ( .A(n4954), .B(n2494), .C(n835), .D(n6781), .Y(n2533) );
  OR3X2 U9844 ( .A(reg_length00[4]), .B(reg_length00[5]), .C(reg_length00[3]), 
        .Y(n2534) );
  OR3X2 U9845 ( .A(n5006), .B(n6987), .C(n7022), .Y(n6988) );
  OR3X2 U9846 ( .A(n7012), .B(n7020), .C(n6988), .Y(n6993) );
  OR4X2 U9847 ( .A(n164), .B(n583), .C(n166), .D(n165), .Y(n6994) );
  OR4X2 U9848 ( .A(n582), .B(n6996), .C(n6995), .D(n6994), .Y(n6997) );
  OR3X2 U9849 ( .A(n878), .B(n7003), .C(n880), .Y(n7005) );
  XNOR2X1 U9850 ( .A(n5377), .B(sub_838_carry_6_), .Y(N5128) );
  XNOR2X1 U9851 ( .A(n5377), .B(sub_844_carry_6_), .Y(N5144) );
  XNOR2X1 U9852 ( .A(n5377), .B(sub_841_carry[6]), .Y(N5136) );
  XOR2X1 U9853 ( .A(n5377), .B(sub_829_carry[6]), .Y(N5104) );
  XOR2X1 U9854 ( .A(n5377), .B(sub_832_carry_6_), .Y(N5112) );
  XNOR2X1 U9855 ( .A(n5378), .B(sub_817_carry_6_), .Y(N5072) );
  XOR2X1 U9856 ( .A(n5377), .B(sub_826_carry_6_), .Y(N5096) );
  XNOR2X1 U9857 ( .A(n5378), .B(N5118), .Y(N5064) );
  XNOR2X1 U9858 ( .A(n5378), .B(sub_820_carry_6_), .Y(N5080) );
  AND2X1 U9859 ( .A(sub_844_carry_5_), .B(n5378), .Y(sub_844_carry_6_) );
  XOR2X1 U9860 ( .A(n5378), .B(sub_844_carry_5_), .Y(N5143) );
  AND2X1 U9861 ( .A(sub_838_carry_5_), .B(n5378), .Y(sub_838_carry_6_) );
  XOR2X1 U9862 ( .A(n5378), .B(sub_838_carry_5_), .Y(N5127) );
  AND2X1 U9863 ( .A(sub_841_carry[5]), .B(n5378), .Y(sub_841_carry[6]) );
  XOR2X1 U9864 ( .A(n5378), .B(sub_841_carry[5]), .Y(N5135) );
  OR2X1 U9865 ( .A(n5378), .B(sub_829_carry[5]), .Y(sub_829_carry[6]) );
  XNOR2X1 U9866 ( .A(sub_829_carry[5]), .B(n5378), .Y(N5103) );
  OR2X1 U9867 ( .A(n5378), .B(sub_826_carry_5_), .Y(sub_826_carry_6_) );
  XNOR2X1 U9868 ( .A(sub_826_carry_5_), .B(n5378), .Y(N5095) );
  OR2X1 U9869 ( .A(n5378), .B(sub_832_carry_5_), .Y(sub_832_carry_6_) );
  XNOR2X1 U9870 ( .A(sub_832_carry_5_), .B(n5378), .Y(N5111) );
  AND2X1 U9871 ( .A(sub_820_carry_5_), .B(N5118), .Y(sub_820_carry_6_) );
  XOR2X1 U9872 ( .A(N5118), .B(sub_820_carry_5_), .Y(N5079) );
  OR2X1 U9873 ( .A(N5118), .B(sub_817_carry_5_), .Y(sub_817_carry_6_) );
  XNOR2X1 U9874 ( .A(sub_817_carry_5_), .B(N5118), .Y(N5071) );
  AND2X1 U9875 ( .A(sub_844_carry_4_), .B(N5118), .Y(sub_844_carry_5_) );
  XOR2X1 U9876 ( .A(N5118), .B(sub_844_carry_4_), .Y(N5142) );
  AND2X1 U9877 ( .A(sub_841_carry[4]), .B(N5118), .Y(sub_841_carry[5]) );
  XOR2X1 U9878 ( .A(N5118), .B(sub_841_carry[4]), .Y(N5134) );
  AND2X1 U9879 ( .A(sub_838_carry_4_), .B(N5118), .Y(sub_838_carry_5_) );
  XOR2X1 U9880 ( .A(N5118), .B(sub_838_carry_4_), .Y(N5126) );
  OR2X1 U9881 ( .A(N5118), .B(sub_832_carry_4_), .Y(sub_832_carry_5_) );
  XNOR2X1 U9882 ( .A(sub_832_carry_4_), .B(N5118), .Y(N5110) );
  OR2X1 U9883 ( .A(N5118), .B(sub_829_carry[4]), .Y(sub_829_carry[5]) );
  XNOR2X1 U9884 ( .A(sub_829_carry[4]), .B(N5118), .Y(N5102) );
  OR2X1 U9885 ( .A(N5118), .B(sub_826_carry_4_), .Y(sub_826_carry_5_) );
  XNOR2X1 U9886 ( .A(sub_826_carry_4_), .B(N5118), .Y(N5094) );
  OR2X1 U9887 ( .A(n5568), .B(sub_820_carry_4_), .Y(sub_820_carry_5_) );
  XNOR2X1 U9888 ( .A(sub_820_carry_4_), .B(n5568), .Y(N5078) );
  AND2X1 U9889 ( .A(sub_817_carry_4_), .B(n5568), .Y(sub_817_carry_5_) );
  XOR2X1 U9890 ( .A(n5568), .B(sub_817_carry_4_), .Y(N5070) );
  AND2X1 U9891 ( .A(sub_844_carry_3_), .B(n5568), .Y(sub_844_carry_4_) );
  XOR2X1 U9892 ( .A(n5568), .B(sub_844_carry_3_), .Y(N5141) );
  AND2X1 U9893 ( .A(sub_841_carry[3]), .B(n5568), .Y(sub_841_carry[4]) );
  XOR2X1 U9894 ( .A(n5568), .B(sub_841_carry[3]), .Y(N5133) );
  AND2X1 U9895 ( .A(sub_838_carry_3_), .B(n5568), .Y(sub_838_carry_4_) );
  XOR2X1 U9896 ( .A(n5568), .B(sub_838_carry_3_), .Y(N5125) );
  OR2X1 U9897 ( .A(n5568), .B(sub_832_carry_3_), .Y(sub_832_carry_4_) );
  XNOR2X1 U9898 ( .A(sub_832_carry_3_), .B(n5568), .Y(N5109) );
  OR2X1 U9899 ( .A(n5568), .B(sub_829_carry[3]), .Y(sub_829_carry[4]) );
  XNOR2X1 U9900 ( .A(sub_829_carry[3]), .B(n5568), .Y(N5101) );
  OR2X1 U9901 ( .A(n5568), .B(sub_826_carry_3_), .Y(sub_826_carry_4_) );
  XNOR2X1 U9902 ( .A(sub_826_carry_3_), .B(n5568), .Y(N5093) );
  OR2X1 U9903 ( .A(N5061), .B(sub_820_carry_3_), .Y(sub_820_carry_4_) );
  XNOR2X1 U9904 ( .A(sub_820_carry_3_), .B(N5061), .Y(N5077) );
  AND2X1 U9905 ( .A(sub_817_carry_3_), .B(N5061), .Y(sub_817_carry_4_) );
  XOR2X1 U9906 ( .A(N5061), .B(sub_817_carry_3_), .Y(N5069) );
  AND2X1 U9907 ( .A(sub_817_carry_2_), .B(n5571), .Y(sub_817_carry_3_) );
  XOR2X1 U9908 ( .A(n5571), .B(sub_817_carry_2_), .Y(N5068) );
  OR2X1 U9909 ( .A(N5061), .B(sub_826_carry_2_), .Y(sub_826_carry_3_) );
  XNOR2X1 U9910 ( .A(sub_826_carry_2_), .B(N5061), .Y(N5092) );
  OR2X1 U9911 ( .A(n5571), .B(sub_820_carry_2_), .Y(sub_820_carry_3_) );
  XNOR2X1 U9912 ( .A(sub_820_carry_2_), .B(n5571), .Y(N5076) );
  AND2X1 U9913 ( .A(sub_838_carry_2_), .B(N5061), .Y(sub_838_carry_3_) );
  XOR2X1 U9914 ( .A(N5061), .B(sub_838_carry_2_), .Y(N5124) );
  AND2X1 U9915 ( .A(sub_844_carry_2_), .B(N5061), .Y(sub_844_carry_3_) );
  XOR2X1 U9916 ( .A(N5061), .B(sub_844_carry_2_), .Y(N5140) );
  AND2X1 U9917 ( .A(n5571), .B(N5061), .Y(sub_841_carry[3]) );
  XOR2X1 U9918 ( .A(N5061), .B(n5571), .Y(N5132) );
  OR2X1 U9919 ( .A(N5061), .B(n5571), .Y(sub_829_carry[3]) );
  XNOR2X1 U9920 ( .A(n5571), .B(N5061), .Y(N5100) );
  OR2X1 U9921 ( .A(N5061), .B(sub_832_carry_2_), .Y(sub_832_carry_3_) );
  XNOR2X1 U9922 ( .A(sub_832_carry_2_), .B(N5061), .Y(N5108) );
  OR2X1 U9923 ( .A(N5059), .B(n5379), .Y(sub_820_carry_2_) );
  XNOR2X1 U9924 ( .A(n5379), .B(N5059), .Y(N5075) );
  AND2X1 U9925 ( .A(n5379), .B(N5059), .Y(sub_817_carry_2_) );
  XOR2X1 U9926 ( .A(N5059), .B(n5379), .Y(N5067) );
  OR2X1 U9927 ( .A(n5571), .B(N5059), .Y(sub_844_carry_2_) );
  XNOR2X1 U9928 ( .A(N5059), .B(n5571), .Y(N5139) );
  AND2X1 U9929 ( .A(N5059), .B(n5571), .Y(sub_838_carry_2_) );
  XOR2X1 U9930 ( .A(n5571), .B(N5059), .Y(N5123) );
  OR2X1 U9931 ( .A(n5571), .B(N5059), .Y(sub_832_carry_2_) );
  XNOR2X1 U9932 ( .A(N5059), .B(n5571), .Y(N5107) );
  AND2X1 U9933 ( .A(N5059), .B(n5571), .Y(sub_826_carry_2_) );
  XOR2X1 U9934 ( .A(n5571), .B(N5059), .Y(N5091) );
  XOR2X1 U9935 ( .A(r889_carry[5]), .B(count_state_idle[5]), .Y(N4526) );
  CLKINVX1 U9936 ( .A(reg_length1[0]), .Y(N7475) );
  OR2X1 U9937 ( .A(reg_length1[1]), .B(reg_length1[0]), .Y(n7048) );
  OAI2BB1X1 U9938 ( .A0N(reg_length1[1]), .A1N(reg_length1[0]), .B0(n7048), 
        .Y(N7476) );
  OR2X1 U9939 ( .A(n7048), .B(reg_length1[2]), .Y(n7049) );
  OAI2BB1X1 U9940 ( .A0N(n7048), .A1N(reg_length1[2]), .B0(n7049), .Y(N7477)
         );
  NOR2X1 U9941 ( .A(n7049), .B(reg_length1[3]), .Y(n7050) );
  OAI2BB1X1 U9942 ( .A0N(n7049), .A1N(reg_length1[3]), .B0(n7052), .Y(N7478)
         );
  XOR2X1 U9943 ( .A(reg_length1[4]), .B(n7050), .Y(N7479) );
  NOR2X1 U9944 ( .A(reg_length1[4]), .B(n7052), .Y(n7051) );
  XOR2X1 U9945 ( .A(reg_length1[5]), .B(n7051), .Y(N7480) );
  CLKINVX1 U9946 ( .A(reg_length2[0]), .Y(N7521) );
  OR2X1 U9947 ( .A(reg_length2[1]), .B(reg_length2[0]), .Y(n7053) );
  OAI2BB1X1 U9948 ( .A0N(reg_length2[1]), .A1N(reg_length2[0]), .B0(n7053), 
        .Y(N7522) );
  OR2X1 U9949 ( .A(n7053), .B(reg_length2[2]), .Y(n7054) );
  OAI2BB1X1 U9950 ( .A0N(n7053), .A1N(reg_length2[2]), .B0(n7054), .Y(N7523)
         );
  NOR2X1 U9951 ( .A(n7054), .B(reg_length2[3]), .Y(n7055) );
  OAI2BB1X1 U9952 ( .A0N(n7054), .A1N(reg_length2[3]), .B0(n7057), .Y(N7524)
         );
  XOR2X1 U9953 ( .A(reg_length2[4]), .B(n7055), .Y(N7525) );
  NOR2X1 U9954 ( .A(reg_length2[4]), .B(n7057), .Y(n7056) );
  XOR2X1 U9955 ( .A(reg_length2[5]), .B(n7056), .Y(N7526) );
  CLKINVX1 U9956 ( .A(reg_length3[0]), .Y(N7565) );
  OR2X1 U9957 ( .A(reg_length3[1]), .B(reg_length3[0]), .Y(n7058) );
  OAI2BB1X1 U9958 ( .A0N(reg_length3[1]), .A1N(reg_length3[0]), .B0(n7058), 
        .Y(N7566) );
  OR2X1 U9959 ( .A(n7058), .B(reg_length3[2]), .Y(n7059) );
  OAI2BB1X1 U9960 ( .A0N(n7058), .A1N(reg_length3[2]), .B0(n7059), .Y(N7567)
         );
  NOR2X1 U9961 ( .A(n7059), .B(reg_length3[3]), .Y(n7060) );
  OAI2BB1X1 U9962 ( .A0N(n7059), .A1N(reg_length3[3]), .B0(n7062), .Y(N7568)
         );
  XOR2X1 U9963 ( .A(reg_length3[4]), .B(n7060), .Y(N7569) );
  NOR2X1 U9964 ( .A(reg_length3[4]), .B(n7062), .Y(n7061) );
  XOR2X1 U9965 ( .A(reg_length3[5]), .B(n7061), .Y(N7570) );
  CLKINVX1 U9966 ( .A(reg_length4[0]), .Y(N7606) );
  OR2X1 U9967 ( .A(reg_length4[1]), .B(reg_length4[0]), .Y(n7063) );
  OAI2BB1X1 U9968 ( .A0N(reg_length4[1]), .A1N(reg_length4[0]), .B0(n7063), 
        .Y(N7607) );
  OR2X1 U9969 ( .A(n7063), .B(reg_length4[2]), .Y(n7064) );
  OAI2BB1X1 U9970 ( .A0N(n7063), .A1N(reg_length4[2]), .B0(n7064), .Y(N7608)
         );
  NOR2X1 U9971 ( .A(n7064), .B(reg_length4[3]), .Y(n7065) );
  OAI2BB1X1 U9972 ( .A0N(n7064), .A1N(reg_length4[3]), .B0(n7067), .Y(N7609)
         );
  XOR2X1 U9973 ( .A(reg_length4[4]), .B(n7065), .Y(N7610) );
  NOR2X1 U9974 ( .A(reg_length4[4]), .B(n7067), .Y(n7066) );
  XOR2X1 U9975 ( .A(reg_length4[5]), .B(n7066), .Y(N7611) );
  OR2X1 U9976 ( .A(reg_length5[1]), .B(reg_length5[0]), .Y(n7068) );
  OAI2BB1X1 U9977 ( .A0N(reg_length5[1]), .A1N(reg_length5[0]), .B0(n7068), 
        .Y(N7648) );
  OR2X1 U9978 ( .A(n7068), .B(reg_length5[2]), .Y(n7069) );
  OAI2BB1X1 U9979 ( .A0N(n7068), .A1N(reg_length5[2]), .B0(n7069), .Y(N7649)
         );
  NOR2X1 U9980 ( .A(n7069), .B(reg_length5[3]), .Y(n7070) );
  OAI2BB1X1 U9981 ( .A0N(n7069), .A1N(reg_length5[3]), .B0(n7072), .Y(N7650)
         );
  XOR2X1 U9982 ( .A(reg_length5[4]), .B(n7070), .Y(N7651) );
  NOR2X1 U9983 ( .A(reg_length5[4]), .B(n7072), .Y(n7071) );
  XOR2X1 U9984 ( .A(reg_length5[5]), .B(n7071), .Y(N7652) );
  CLKINVX1 U9985 ( .A(reg_length6[0]), .Y(N7688) );
  OR2X1 U9986 ( .A(reg_length6[1]), .B(reg_length6[0]), .Y(n7073) );
  OAI2BB1X1 U9987 ( .A0N(reg_length6[1]), .A1N(reg_length6[0]), .B0(n7073), 
        .Y(N7689) );
  OR2X1 U9988 ( .A(n7073), .B(reg_length6[2]), .Y(n7074) );
  OAI2BB1X1 U9989 ( .A0N(n7073), .A1N(reg_length6[2]), .B0(n7074), .Y(N7690)
         );
  NOR2X1 U9990 ( .A(n7074), .B(reg_length6[3]), .Y(n7075) );
  OAI2BB1X1 U9991 ( .A0N(n7074), .A1N(reg_length6[3]), .B0(n7077), .Y(N7691)
         );
  XOR2X1 U9992 ( .A(reg_length6[4]), .B(n7075), .Y(N7692) );
  NOR2X1 U9993 ( .A(reg_length6[4]), .B(n7077), .Y(n7076) );
  XOR2X1 U9994 ( .A(reg_length6[5]), .B(n7076), .Y(N7693) );
  CLKINVX1 U9995 ( .A(reg_length7[0]), .Y(N7727) );
  OR2X1 U9996 ( .A(reg_length7[1]), .B(reg_length7[0]), .Y(n7078) );
  OAI2BB1X1 U9997 ( .A0N(reg_length7[1]), .A1N(reg_length7[0]), .B0(n7078), 
        .Y(N7728) );
  OR2X1 U9998 ( .A(n7078), .B(reg_length7[2]), .Y(n7079) );
  OAI2BB1X1 U9999 ( .A0N(n7078), .A1N(reg_length7[2]), .B0(n7079), .Y(N7729)
         );
  NOR2X1 U10000 ( .A(n7079), .B(reg_length7[3]), .Y(n7080) );
  OAI2BB1X1 U10001 ( .A0N(n7079), .A1N(reg_length7[3]), .B0(n7082), .Y(N7730)
         );
  XOR2X1 U10002 ( .A(reg_length7[4]), .B(n7080), .Y(N7731) );
  NOR2X1 U10003 ( .A(reg_length7[4]), .B(n7082), .Y(n7081) );
  OR2X1 U10004 ( .A(reg_length8[1]), .B(reg_length8[0]), .Y(n7083) );
  OAI2BB1X1 U10005 ( .A0N(reg_length8[1]), .A1N(reg_length8[0]), .B0(n7083), 
        .Y(N7764) );
  OR2X1 U10006 ( .A(n7083), .B(reg_length8[2]), .Y(n7084) );
  OAI2BB1X1 U10007 ( .A0N(n7083), .A1N(reg_length8[2]), .B0(n7084), .Y(N7765)
         );
  NOR2X1 U10008 ( .A(n7084), .B(reg_length8[3]), .Y(n7085) );
  OAI2BB1X1 U10009 ( .A0N(n7084), .A1N(reg_length8[3]), .B0(n7086), .Y(N7766)
         );
  XOR2X1 U10010 ( .A(reg_length8[4]), .B(n7085), .Y(N7767) );
  CLKINVX1 U10011 ( .A(reg_length9[0]), .Y(N7799) );
  OR2X1 U10012 ( .A(reg_length9[1]), .B(reg_length9[0]), .Y(n7087) );
  OAI2BB1X1 U10013 ( .A0N(reg_length9[1]), .A1N(reg_length9[0]), .B0(n7087), 
        .Y(N7800) );
  OR2X1 U10014 ( .A(n7087), .B(reg_length9[2]), .Y(n7088) );
  OAI2BB1X1 U10015 ( .A0N(n7087), .A1N(reg_length9[2]), .B0(n7088), .Y(N7801)
         );
  NOR2X1 U10016 ( .A(n7088), .B(reg_length9[3]), .Y(n7089) );
  OAI2BB1X1 U10017 ( .A0N(n7088), .A1N(reg_length9[3]), .B0(n7090), .Y(N7802)
         );
  XOR2X1 U10018 ( .A(reg_length9[4]), .B(n7089), .Y(N7803) );
  CLKINVX1 U10019 ( .A(n5364), .Y(N7835) );
  OR2X1 U10020 ( .A(reg_length10[1]), .B(n5364), .Y(n7091) );
  OAI2BB1X1 U10021 ( .A0N(reg_length10[1]), .A1N(n5364), .B0(n7091), .Y(N7836)
         );
  OR2X1 U10022 ( .A(n7091), .B(reg_length10[2]), .Y(n7092) );
  OAI2BB1X1 U10023 ( .A0N(n7091), .A1N(reg_length10[2]), .B0(n7092), .Y(N7837)
         );
  NOR2X1 U10024 ( .A(n7092), .B(reg_length10[3]), .Y(n7093) );
  OAI2BB1X1 U10025 ( .A0N(n7092), .A1N(reg_length10[3]), .B0(n7095), .Y(N7838)
         );
  XOR2X1 U10026 ( .A(reg_length10[4]), .B(n7093), .Y(N7839) );
  NOR2X1 U10027 ( .A(reg_length10[4]), .B(n7095), .Y(n7094) );
  XOR2X1 U10028 ( .A(reg_length10[5]), .B(n7094), .Y(N7840) );
  CLKINVX1 U10029 ( .A(reg_length11[0]), .Y(N7871) );
  OR2X1 U10030 ( .A(reg_length11[1]), .B(reg_length11[0]), .Y(n7096) );
  OAI2BB1X1 U10031 ( .A0N(reg_length11[1]), .A1N(reg_length11[0]), .B0(n7096), 
        .Y(N7872) );
  OR2X1 U10032 ( .A(n7096), .B(reg_length11[2]), .Y(n7097) );
  OAI2BB1X1 U10033 ( .A0N(n7096), .A1N(reg_length11[2]), .B0(n7097), .Y(N7873)
         );
  NOR2X1 U10034 ( .A(n7097), .B(reg_length11[3]), .Y(n7098) );
  OAI2BB1X1 U10035 ( .A0N(n7097), .A1N(reg_length11[3]), .B0(n7099), .Y(N7874)
         );
  XOR2X1 U10036 ( .A(reg_length11[4]), .B(n7098), .Y(N7875) );
  CLKINVX1 U10037 ( .A(n5365), .Y(N7907) );
  OR2X1 U10038 ( .A(reg_length12[1]), .B(n5365), .Y(n7100) );
  OAI2BB1X1 U10039 ( .A0N(reg_length12[1]), .A1N(n5365), .B0(n7100), .Y(N7908)
         );
  OR2X1 U10040 ( .A(n7100), .B(reg_length12[2]), .Y(n7101) );
  OAI2BB1X1 U10041 ( .A0N(n7100), .A1N(reg_length12[2]), .B0(n7101), .Y(N7909)
         );
  NOR2X1 U10042 ( .A(n7101), .B(reg_length12[3]), .Y(n7102) );
  OAI2BB1X1 U10043 ( .A0N(n7101), .A1N(reg_length12[3]), .B0(n7103), .Y(N7910)
         );
  XOR2X1 U10044 ( .A(reg_length12[4]), .B(n7102), .Y(N7911) );
  CLKINVX1 U10045 ( .A(reg_length13[0]), .Y(N7943) );
  OR2X1 U10046 ( .A(reg_length13[1]), .B(reg_length13[0]), .Y(n7104) );
  OAI2BB1X1 U10047 ( .A0N(reg_length13[1]), .A1N(reg_length13[0]), .B0(n7104), 
        .Y(N7944) );
  OR2X1 U10048 ( .A(n7104), .B(reg_length13[2]), .Y(n7105) );
  OAI2BB1X1 U10049 ( .A0N(n7104), .A1N(reg_length13[2]), .B0(n7105), .Y(N7945)
         );
  NOR2X1 U10050 ( .A(n7105), .B(reg_length13[3]), .Y(n7106) );
  OAI2BB1X1 U10051 ( .A0N(n7105), .A1N(reg_length13[3]), .B0(n7107), .Y(N7946)
         );
  XOR2X1 U10052 ( .A(reg_length13[4]), .B(n7106), .Y(N7947) );
  OR2X1 U10053 ( .A(reg_length14[1]), .B(reg_length14[0]), .Y(n7108) );
  OAI2BB1X1 U10054 ( .A0N(reg_length14[1]), .A1N(reg_length14[0]), .B0(n7108), 
        .Y(N7980) );
  OR2X1 U10055 ( .A(n7108), .B(reg_length14[2]), .Y(n7109) );
  OAI2BB1X1 U10056 ( .A0N(n7108), .A1N(reg_length14[2]), .B0(n7109), .Y(N7981)
         );
  NOR2X1 U10057 ( .A(n7109), .B(reg_length14[3]), .Y(n7110) );
  OAI2BB1X1 U10058 ( .A0N(n7109), .A1N(reg_length14[3]), .B0(n7111), .Y(N7982)
         );
  XOR2X1 U10059 ( .A(reg_length14[4]), .B(n7110), .Y(N7983) );
  NOR4X1 U10060 ( .A(N5059), .B(n5379), .C(n5380), .D(count[3]), .Y(n7112) );
  NOR4BX1 U10061 ( .AN(n7112), .B(count[2]), .C(count[0]), .D(count[1]), .Y(
        n7113) );
  NAND4BX1 U10062 ( .AN(n7113), .B(n5571), .C(n5568), .D(N5061), .Y(N5018) );
  OR4X1 U10063 ( .A(n5379), .B(n5380), .C(n5571), .D(N5059), .Y(n7115) );
  OR4X1 U10064 ( .A(count[1]), .B(count[0]), .C(count[3]), .D(count[2]), .Y(
        n7114) );
  OAI211X1 U10065 ( .A0(n7115), .A1(n7114), .B0(N5061), .C0(n5568), .Y(N5016)
         );
  OR4X1 U10066 ( .A(n5380), .B(count[3]), .C(N5059), .D(n5379), .Y(n7116) );
  OR4X1 U10067 ( .A(count[2]), .B(count[1]), .C(count[0]), .D(n7116), .Y(n7117) );
  AOI32X1 U10068 ( .A0(n5571), .A1(n7117), .A2(n5568), .B0(N5061), .B1(n5568), 
        .Y(N5014) );
  NOR4X1 U10069 ( .A(count[3]), .B(count[2]), .C(count[1]), .D(count[0]), .Y(
        n7120) );
  NOR2X1 U10070 ( .A(N5061), .B(n5571), .Y(n7118) );
  NOR4BX1 U10071 ( .AN(n7118), .B(n5379), .C(n5380), .D(N5059), .Y(n7119) );
  OAI2BB1X1 U10072 ( .A0N(n7120), .A1N(n7119), .B0(n5568), .Y(N5012) );
  NOR4X1 U10073 ( .A(count[3]), .B(count[2]), .C(count[1]), .D(count[0]), .Y(
        n7123) );
  NOR4X1 U10074 ( .A(n5568), .B(N5059), .C(n5379), .D(n5380), .Y(n7122) );
  AOI21X1 U10075 ( .A0(N5061), .A1(n5571), .B0(n5568), .Y(n7121) );
  OAI2BB1X1 U10076 ( .A0N(n7123), .A1N(n7122), .B0(n7124), .Y(N5010) );
  NOR4X1 U10077 ( .A(count[3]), .B(count[2]), .C(count[1]), .D(count[0]), .Y(
        n7126) );
  NOR4X1 U10078 ( .A(n5571), .B(N5059), .C(n5379), .D(n5380), .Y(n7125) );
  NAND2X1 U10079 ( .A(n7126), .B(n7125), .Y(n7127) );
  AOI21X1 U10080 ( .A0(N5061), .A1(n7127), .B0(n5568), .Y(N5008) );
  OR4X1 U10081 ( .A(n5380), .B(count[3]), .C(N5059), .D(n5379), .Y(n7128) );
  OR4X1 U10082 ( .A(count[2]), .B(count[1]), .C(count[0]), .D(n7128), .Y(n7129) );
  AOI211X1 U10083 ( .A0(n5571), .A1(n7129), .B0(n5568), .C0(N5061), .Y(N5006)
         );
  AOI211X1 U10084 ( .A0(n5374), .A1(n5375), .B0(n5373), .C0(reg_invalid2[4]), 
        .Y(n7130) );
  NOR4BX1 U10085 ( .AN(n7130), .B(reg_invalid2[8]), .C(reg_invalid2[6]), .D(
        reg_invalid2[7]), .Y(N8480) );
  AOI211X1 U10086 ( .A0(n5374), .A1(n5375), .B0(n5373), .C0(reg_invalid2[4]), 
        .Y(n7132) );
  NOR3X1 U10087 ( .A(reg_invalid2[6]), .B(reg_invalid2[8]), .C(reg_invalid2[7]), .Y(n7131) );
  NAND2X1 U10088 ( .A(n7132), .B(n7131), .Y(N7419) );
  OR2X1 U10089 ( .A(reg_invalid2[8]), .B(reg_invalid2[7]), .Y(n7133) );
  AOI21X1 U10090 ( .A0(reg_invalid2[6]), .A1(n5373), .B0(n7133), .Y(n7135) );
  OAI211X1 U10091 ( .A0(n5375), .A1(n5376), .B0(n5374), .C0(reg_invalid2[4]), 
        .Y(n7134) );
  AOI22X1 U10092 ( .A0(n7135), .A1(n7331), .B0(n7135), .B1(n7134), .Y(N4685)
         );
endmodule


module MMSA_DW01_add_44 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n63, n64, n65, n66, n67, n68, n69, n70, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n128, n129, n130, n131, n132, n133,
         n136, n137, n138, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n153, n155, n156, n157, n158, n160, n163,
         n164, n165, n166, n167, n169, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n201, n203, n204, n205, n206, n207, n209, n211, n212, n213,
         n214, n215, n217, n219, n220, n221, n222, n223, n225, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n237, n239, n240, n241,
         n242, n243, n245, n247, n253, n254, n255, n256, n270, n273, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435;

  AOI21X1 U17 ( .A0(n51), .A1(n68), .B0(n52), .Y(n50) );
  AOI21X1 U27 ( .A0(n58), .A1(n86), .B0(n59), .Y(n57) );
  AOI21X1 U39 ( .A0(n86), .A1(n67), .B0(n68), .Y(n66) );
  AOI21X1 U53 ( .A0(n86), .A1(n78), .B0(n79), .Y(n77) );
  AOI21X1 U77 ( .A0(n104), .A1(n96), .B0(n97), .Y(n95) );
  AOI21X1 U108 ( .A0(n131), .A1(n118), .B0(n119), .Y(n117) );
  AOI21X1 U116 ( .A0(n123), .A1(n143), .B0(n124), .Y(n122) );
  AOI21X1 U126 ( .A0(n143), .A1(n130), .B0(n131), .Y(n129) );
  AOI21X1 U138 ( .A0(n143), .A1(n270), .B0(n140), .Y(n138) );
  AOI21X1 U157 ( .A0(n430), .A1(n160), .B0(n153), .Y(n151) );
  NOR2X2 U222 ( .A(B[16]), .B(A[16]), .Y(n190) );
  NOR2X2 U228 ( .A(B[15]), .B(A[15]), .Y(n193) );
  OAI21X1 U340 ( .A0(n165), .A1(n167), .B0(n166), .Y(n164) );
  AOI21X1 U341 ( .A0(n145), .A1(n164), .B0(n146), .Y(n144) );
  NOR2X1 U342 ( .A(B[18]), .B(A[18]), .Y(n181) );
  NOR2X1 U343 ( .A(n112), .B(n109), .Y(n103) );
  NOR2X1 U344 ( .A(n80), .B(n73), .Y(n67) );
  OAI21X1 U345 ( .A0(n116), .A1(n144), .B0(n117), .Y(n115) );
  NAND2X1 U346 ( .A(n130), .B(n118), .Y(n116) );
  AOI21X1 U347 ( .A0(n172), .A1(n427), .B0(n169), .Y(n167) );
  NOR2X1 U348 ( .A(B[30]), .B(A[30]), .Y(n112) );
  OAI21X1 U349 ( .A0(n173), .A1(n175), .B0(n174), .Y(n172) );
  NOR2X1 U350 ( .A(B[28]), .B(A[28]), .Y(n125) );
  NOR2X1 U351 ( .A(n423), .B(n189), .Y(n187) );
  OAI21X1 U352 ( .A0(n190), .A1(n194), .B0(n191), .Y(n189) );
  AND2X1 U353 ( .A(n188), .B(n196), .Y(n423) );
  NOR2X1 U354 ( .A(B[27]), .B(A[27]), .Y(n136) );
  NOR2X1 U355 ( .A(B[29]), .B(A[29]), .Y(n120) );
  OAI21X2 U356 ( .A0(n187), .A1(n185), .B0(n186), .Y(n184) );
  NAND2XL U357 ( .A(n85), .B(n67), .Y(n65) );
  CLKINVXL U358 ( .A(n81), .Y(n79) );
  NOR2X1 U359 ( .A(B[33]), .B(A[33]), .Y(n91) );
  OAI21XL U360 ( .A0(n114), .A1(n65), .B0(n66), .Y(n64) );
  OAI21XL U361 ( .A0(n114), .A1(n101), .B0(n102), .Y(n100) );
  OAI21XL U362 ( .A0(n114), .A1(n56), .B0(n57), .Y(n55) );
  OAI21XL U363 ( .A0(n114), .A1(n76), .B0(n77), .Y(n75) );
  OAI21X1 U364 ( .A0(n73), .A1(n81), .B0(n74), .Y(n68) );
  OAI21X1 U365 ( .A0(n233), .A1(n235), .B0(n234), .Y(n232) );
  INVX1 U366 ( .A(n84), .Y(n86) );
  INVX2 U367 ( .A(n115), .Y(n114) );
  CLKINVXL U368 ( .A(n104), .Y(n102) );
  CLKINVXL U369 ( .A(n103), .Y(n101) );
  OAI21XL U370 ( .A0(n114), .A1(n83), .B0(n84), .Y(n82) );
  NAND2XL U371 ( .A(n89), .B(n103), .Y(n83) );
  CLKINVXL U372 ( .A(n144), .Y(n143) );
  OAI21XL U373 ( .A0(n163), .A1(n150), .B0(n151), .Y(n149) );
  CLKINVXL U374 ( .A(n130), .Y(n132) );
  CLKINVXL U375 ( .A(n184), .Y(n183) );
  CLKINVXL U376 ( .A(n196), .Y(n195) );
  OAI21X1 U377 ( .A0(n142), .A1(n136), .B0(n137), .Y(n131) );
  CLKINVXL U378 ( .A(n99), .Y(n97) );
  CLKINVXL U379 ( .A(n98), .Y(n96) );
  CLKINVX2 U380 ( .A(n157), .Y(n273) );
  NAND2XL U381 ( .A(n96), .B(n99), .Y(n8) );
  OAI21XL U382 ( .A0(n163), .A1(n157), .B0(n158), .Y(n156) );
  OAI21XL U383 ( .A0(n53), .A1(n63), .B0(n54), .Y(n52) );
  INVX1 U384 ( .A(n232), .Y(n231) );
  CLKINVXL U385 ( .A(n141), .Y(n270) );
  CLKINVXL U386 ( .A(n80), .Y(n78) );
  NAND2BXL U387 ( .AN(n125), .B(n128), .Y(n12) );
  NAND2BXL U388 ( .AN(n91), .B(n92), .Y(n7) );
  NAND2XL U389 ( .A(n273), .B(n158), .Y(n17) );
  NAND2BXL U390 ( .AN(n185), .B(n186), .Y(n23) );
  NAND2BXL U391 ( .AN(n190), .B(n191), .Y(n24) );
  NAND2XL U392 ( .A(n429), .B(n211), .Y(n29) );
  NAND2XL U393 ( .A(n432), .B(n219), .Y(n31) );
  OR2XL U394 ( .A(B[24]), .B(A[24]), .Y(n430) );
  NAND2XL U395 ( .A(B[24]), .B(A[24]), .Y(n155) );
  NAND2XL U396 ( .A(B[26]), .B(A[26]), .Y(n142) );
  NAND2XL U397 ( .A(B[23]), .B(A[23]), .Y(n158) );
  NAND2XL U398 ( .A(B[30]), .B(A[30]), .Y(n113) );
  NAND2XL U399 ( .A(B[18]), .B(A[18]), .Y(n182) );
  NAND2XL U400 ( .A(B[15]), .B(A[15]), .Y(n194) );
  NAND2XL U401 ( .A(B[8]), .B(A[8]), .Y(n222) );
  OR2XL U402 ( .A(B[13]), .B(A[13]), .Y(n425) );
  NAND2XL U403 ( .A(B[13]), .B(A[13]), .Y(n203) );
  OR2XL U404 ( .A(B[21]), .B(A[21]), .Y(n427) );
  OR2XL U405 ( .A(B[7]), .B(A[7]), .Y(n428) );
  NAND2XL U406 ( .A(B[21]), .B(A[21]), .Y(n171) );
  NAND2XL U407 ( .A(B[11]), .B(A[11]), .Y(n211) );
  NAND2XL U408 ( .A(B[7]), .B(A[7]), .Y(n227) );
  NAND2XL U409 ( .A(B[14]), .B(A[14]), .Y(n198) );
  NAND2XL U410 ( .A(B[10]), .B(A[10]), .Y(n214) );
  NAND2XL U411 ( .A(B[34]), .B(A[34]), .Y(n81) );
  NAND2XL U412 ( .A(B[22]), .B(A[22]), .Y(n166) );
  NAND2XL U413 ( .A(B[36]), .B(A[36]), .Y(n63) );
  OR2XL U414 ( .A(B[4]), .B(A[4]), .Y(n426) );
  NAND2XL U415 ( .A(B[4]), .B(A[4]), .Y(n239) );
  NAND2XL U416 ( .A(n434), .B(A[38]), .Y(n45) );
  NAND2BX1 U417 ( .AN(n41), .B(n42), .Y(n1) );
  INVX2 U418 ( .A(n435), .Y(n434) );
  INVX2 U419 ( .A(B[38]), .Y(n435) );
  INVX2 U420 ( .A(n83), .Y(n85) );
  AOI21X1 U421 ( .A0(n115), .A1(n47), .B0(n48), .Y(n46) );
  OAI21X1 U422 ( .A0(n84), .A1(n49), .B0(n50), .Y(n48) );
  NOR2X1 U423 ( .A(n49), .B(n83), .Y(n47) );
  NAND2X1 U424 ( .A(n67), .B(n51), .Y(n49) );
  INVX2 U425 ( .A(n67), .Y(n69) );
  CLKINVXL U426 ( .A(n164), .Y(n163) );
  NOR2X1 U427 ( .A(n60), .B(n53), .Y(n51) );
  OAI21X1 U428 ( .A0(n46), .A1(n44), .B0(n45), .Y(n43) );
  NAND2XL U429 ( .A(n58), .B(n85), .Y(n56) );
  NOR2X1 U430 ( .A(n69), .B(n60), .Y(n58) );
  OAI21X1 U431 ( .A0(n70), .A1(n60), .B0(n63), .Y(n59) );
  CLKINVXL U432 ( .A(n68), .Y(n70) );
  NOR2X1 U433 ( .A(n141), .B(n136), .Y(n130) );
  OAI21XL U434 ( .A0(n120), .A1(n128), .B0(n121), .Y(n119) );
  OAI21XL U435 ( .A0(n114), .A1(n112), .B0(n113), .Y(n111) );
  OAI21XL U436 ( .A0(n114), .A1(n94), .B0(n95), .Y(n93) );
  NAND2XL U437 ( .A(n103), .B(n96), .Y(n94) );
  NAND2XL U438 ( .A(n85), .B(n78), .Y(n76) );
  NOR2X1 U439 ( .A(n125), .B(n120), .Y(n118) );
  AOI21X1 U440 ( .A0(n176), .A1(n184), .B0(n177), .Y(n175) );
  OAI21X1 U441 ( .A0(n178), .A1(n182), .B0(n179), .Y(n177) );
  NOR2X1 U442 ( .A(n181), .B(n178), .Y(n176) );
  INVX2 U443 ( .A(n171), .Y(n169) );
  OAI21X1 U444 ( .A0(n151), .A1(n147), .B0(n148), .Y(n146) );
  NOR2X1 U445 ( .A(n150), .B(n147), .Y(n145) );
  NOR2X1 U446 ( .A(n193), .B(n190), .Y(n188) );
  OAI21XL U447 ( .A0(n133), .A1(n125), .B0(n128), .Y(n124) );
  NOR2X1 U448 ( .A(n132), .B(n125), .Y(n123) );
  CLKINVXL U449 ( .A(n131), .Y(n133) );
  OAI21X1 U450 ( .A0(n199), .A1(n197), .B0(n198), .Y(n196) );
  INVX2 U451 ( .A(n142), .Y(n140) );
  AOI21X1 U452 ( .A0(n204), .A1(n425), .B0(n201), .Y(n199) );
  INVX2 U453 ( .A(n203), .Y(n201) );
  AOI21X1 U454 ( .A0(n429), .A1(n212), .B0(n209), .Y(n207) );
  INVX2 U455 ( .A(n211), .Y(n209) );
  AOI21X1 U456 ( .A0(n426), .A1(n240), .B0(n237), .Y(n235) );
  INVX2 U457 ( .A(n239), .Y(n237) );
  AOI21X1 U458 ( .A0(n228), .A1(n428), .B0(n225), .Y(n223) );
  INVX2 U459 ( .A(n227), .Y(n225) );
  AOI21X1 U460 ( .A0(n220), .A1(n432), .B0(n217), .Y(n215) );
  INVX2 U461 ( .A(n219), .Y(n217) );
  OAI21X1 U462 ( .A0(n221), .A1(n223), .B0(n222), .Y(n220) );
  OAI21X1 U463 ( .A0(n205), .A1(n207), .B0(n206), .Y(n204) );
  OAI21X1 U464 ( .A0(n229), .A1(n231), .B0(n230), .Y(n228) );
  OAI21X1 U465 ( .A0(n213), .A1(n215), .B0(n214), .Y(n212) );
  INVX2 U466 ( .A(n155), .Y(n153) );
  INVX2 U467 ( .A(n158), .Y(n160) );
  AOI21X1 U468 ( .A0(n89), .A1(n104), .B0(n90), .Y(n84) );
  OAI21X1 U469 ( .A0(n91), .A1(n99), .B0(n92), .Y(n90) );
  NOR2X1 U470 ( .A(n91), .B(n98), .Y(n89) );
  AOI21X1 U471 ( .A0(n431), .A1(n424), .B0(n245), .Y(n243) );
  INVX2 U472 ( .A(n247), .Y(n245) );
  OAI21X1 U473 ( .A0(n241), .A1(n243), .B0(n242), .Y(n240) );
  OAI21X1 U474 ( .A0(n109), .A1(n113), .B0(n110), .Y(n104) );
  NAND2BX1 U475 ( .AN(n44), .B(n45), .Y(n2) );
  NAND2X1 U476 ( .A(n273), .B(n430), .Y(n150) );
  OAI2BB1X1 U477 ( .A0N(n433), .A1N(n254), .B0(n253), .Y(n424) );
  NAND2BX1 U478 ( .AN(n53), .B(n54), .Y(n3) );
  NAND2BX1 U479 ( .AN(n60), .B(n63), .Y(n4) );
  NAND2XL U480 ( .A(n78), .B(n81), .Y(n6) );
  NAND2BX1 U481 ( .AN(n73), .B(n74), .Y(n5) );
  NAND2BX1 U482 ( .AN(n136), .B(n137), .Y(n13) );
  NAND2BX1 U483 ( .AN(n120), .B(n121), .Y(n11) );
  NAND2BX1 U484 ( .AN(n112), .B(n113), .Y(n10) );
  NAND2BX1 U485 ( .AN(n147), .B(n148), .Y(n15) );
  NAND2X1 U486 ( .A(n270), .B(n142), .Y(n14) );
  INVX2 U487 ( .A(n256), .Y(n254) );
  NAND2BX1 U488 ( .AN(n109), .B(n110), .Y(n9) );
  NAND2X1 U489 ( .A(n427), .B(n171), .Y(n19) );
  NAND2BX1 U490 ( .AN(n173), .B(n174), .Y(n20) );
  NAND2X1 U491 ( .A(n430), .B(n155), .Y(n16) );
  NAND2BX1 U492 ( .AN(n165), .B(n166), .Y(n18) );
  OAI21XL U493 ( .A0(n183), .A1(n181), .B0(n182), .Y(n180) );
  NAND2BX1 U494 ( .AN(n178), .B(n179), .Y(n21) );
  NAND2BX1 U495 ( .AN(n181), .B(n182), .Y(n22) );
  OAI21XL U496 ( .A0(n195), .A1(n193), .B0(n194), .Y(n192) );
  NAND2BX1 U497 ( .AN(n197), .B(n198), .Y(n26) );
  NAND2BX1 U498 ( .AN(n193), .B(n194), .Y(n25) );
  NAND2X1 U499 ( .A(n425), .B(n203), .Y(n27) );
  NAND2BX1 U500 ( .AN(n205), .B(n206), .Y(n28) );
  NAND2BX1 U501 ( .AN(n213), .B(n214), .Y(n30) );
  NAND2BX1 U502 ( .AN(n221), .B(n222), .Y(n32) );
  NAND2X1 U503 ( .A(n428), .B(n227), .Y(n33) );
  NAND2BX1 U504 ( .AN(n229), .B(n230), .Y(n34) );
  NAND2BX1 U505 ( .AN(n233), .B(n234), .Y(n35) );
  NAND2X1 U506 ( .A(n426), .B(n239), .Y(n36) );
  NAND2BX1 U507 ( .AN(n241), .B(n242), .Y(n37) );
  NAND2X1 U508 ( .A(n431), .B(n247), .Y(n38) );
  NAND2X1 U509 ( .A(n433), .B(n253), .Y(n39) );
  NOR2X1 U510 ( .A(B[37]), .B(A[37]), .Y(n53) );
  XNOR2X1 U511 ( .A(n43), .B(n1), .Y(SUM[39]) );
  NOR2X1 U512 ( .A(B[34]), .B(A[34]), .Y(n80) );
  NOR2X1 U513 ( .A(B[36]), .B(A[36]), .Y(n60) );
  NOR2X1 U514 ( .A(B[35]), .B(A[35]), .Y(n73) );
  XNOR2X1 U515 ( .A(n55), .B(n3), .Y(SUM[37]) );
  XOR2X1 U516 ( .A(n46), .B(n2), .Y(SUM[38]) );
  XNOR2X1 U517 ( .A(n100), .B(n8), .Y(SUM[32]) );
  XNOR2X1 U518 ( .A(n111), .B(n9), .Y(SUM[31]) );
  XNOR2X1 U519 ( .A(n93), .B(n7), .Y(SUM[33]) );
  XNOR2X1 U520 ( .A(n82), .B(n6), .Y(SUM[34]) );
  XNOR2X1 U521 ( .A(n64), .B(n4), .Y(SUM[36]) );
  XNOR2X1 U522 ( .A(n75), .B(n5), .Y(SUM[35]) );
  NAND2XL U523 ( .A(B[35]), .B(A[35]), .Y(n74) );
  NAND2XL U524 ( .A(B[37]), .B(A[37]), .Y(n54) );
  NOR2X1 U525 ( .A(B[19]), .B(A[19]), .Y(n178) );
  XOR2X1 U526 ( .A(n122), .B(n11), .Y(SUM[29]) );
  NOR2X1 U527 ( .A(B[14]), .B(A[14]), .Y(n197) );
  NOR2X1 U528 ( .A(B[31]), .B(A[31]), .Y(n109) );
  XOR2X1 U529 ( .A(n129), .B(n12), .Y(SUM[28]) );
  XOR2X1 U530 ( .A(n138), .B(n13), .Y(SUM[27]) );
  NOR2X1 U531 ( .A(B[20]), .B(A[20]), .Y(n173) );
  NOR2X1 U532 ( .A(B[26]), .B(A[26]), .Y(n141) );
  XOR2X1 U533 ( .A(n114), .B(n10), .Y(SUM[30]) );
  NOR2X1 U534 ( .A(B[17]), .B(A[17]), .Y(n185) );
  NOR2X1 U535 ( .A(B[12]), .B(A[12]), .Y(n205) );
  NOR2X1 U536 ( .A(B[5]), .B(A[5]), .Y(n233) );
  NOR2X1 U537 ( .A(B[6]), .B(A[6]), .Y(n229) );
  NOR2X1 U538 ( .A(B[25]), .B(A[25]), .Y(n147) );
  NOR2X1 U539 ( .A(B[10]), .B(A[10]), .Y(n213) );
  NAND2XL U540 ( .A(B[20]), .B(A[20]), .Y(n174) );
  OR2XL U541 ( .A(B[11]), .B(A[11]), .Y(n429) );
  NAND2XL U542 ( .A(B[19]), .B(A[19]), .Y(n179) );
  NOR2X1 U543 ( .A(B[32]), .B(A[32]), .Y(n98) );
  OR2XL U544 ( .A(B[2]), .B(A[2]), .Y(n431) );
  NAND2XL U545 ( .A(B[27]), .B(A[27]), .Y(n137) );
  NAND2XL U546 ( .A(B[28]), .B(A[28]), .Y(n128) );
  NAND2XL U547 ( .A(B[16]), .B(A[16]), .Y(n191) );
  NOR2X1 U548 ( .A(n434), .B(A[38]), .Y(n44) );
  NOR2X1 U549 ( .A(B[3]), .B(A[3]), .Y(n241) );
  OR2XL U550 ( .A(B[9]), .B(A[9]), .Y(n432) );
  NAND2XL U551 ( .A(B[5]), .B(A[5]), .Y(n234) );
  NAND2XL U552 ( .A(B[12]), .B(A[12]), .Y(n206) );
  NOR2X1 U553 ( .A(B[23]), .B(A[23]), .Y(n157) );
  NAND2XL U554 ( .A(B[29]), .B(A[29]), .Y(n121) );
  NAND2X1 U555 ( .A(B[32]), .B(A[32]), .Y(n99) );
  NAND2XL U556 ( .A(B[17]), .B(A[17]), .Y(n186) );
  NAND2XL U557 ( .A(B[33]), .B(A[33]), .Y(n92) );
  NAND2X1 U558 ( .A(n434), .B(A[39]), .Y(n42) );
  NOR2X1 U559 ( .A(n434), .B(A[39]), .Y(n41) );
  OR2XL U560 ( .A(B[1]), .B(A[1]), .Y(n433) );
  NAND2XL U561 ( .A(B[31]), .B(A[31]), .Y(n110) );
  NAND2XL U562 ( .A(B[6]), .B(A[6]), .Y(n230) );
  NAND2XL U563 ( .A(B[9]), .B(A[9]), .Y(n219) );
  NAND2XL U564 ( .A(B[2]), .B(A[2]), .Y(n247) );
  NOR2X1 U565 ( .A(B[8]), .B(A[8]), .Y(n221) );
  NAND2XL U566 ( .A(B[25]), .B(A[25]), .Y(n148) );
  XNOR2X1 U567 ( .A(n143), .B(n14), .Y(SUM[26]) );
  NAND2XL U568 ( .A(B[1]), .B(A[1]), .Y(n253) );
  NAND2XL U569 ( .A(B[3]), .B(A[3]), .Y(n242) );
  XNOR2X1 U570 ( .A(n156), .B(n16), .Y(SUM[24]) );
  XNOR2X1 U571 ( .A(n149), .B(n15), .Y(SUM[25]) );
  NOR2X1 U572 ( .A(B[22]), .B(A[22]), .Y(n165) );
  XOR2X1 U573 ( .A(n163), .B(n17), .Y(SUM[23]) );
  NAND2X1 U574 ( .A(B[0]), .B(A[0]), .Y(n256) );
  XOR2XL U575 ( .A(n18), .B(n167), .Y(SUM[22]) );
  XNOR2X1 U576 ( .A(n172), .B(n19), .Y(SUM[21]) );
  XOR2XL U577 ( .A(n20), .B(n175), .Y(SUM[20]) );
  XNOR2X1 U578 ( .A(n180), .B(n21), .Y(SUM[19]) );
  XOR2X1 U579 ( .A(n183), .B(n22), .Y(SUM[18]) );
  XOR2X1 U580 ( .A(n187), .B(n23), .Y(SUM[17]) );
  XNOR2X1 U581 ( .A(n192), .B(n24), .Y(SUM[16]) );
  XOR2X1 U582 ( .A(n25), .B(n195), .Y(SUM[15]) );
  XOR2XL U583 ( .A(n26), .B(n199), .Y(SUM[14]) );
  XNOR2XL U584 ( .A(n27), .B(n204), .Y(SUM[13]) );
  XOR2XL U585 ( .A(n28), .B(n207), .Y(SUM[12]) );
  XNOR2XL U586 ( .A(n29), .B(n212), .Y(SUM[11]) );
  XOR2XL U587 ( .A(n30), .B(n215), .Y(SUM[10]) );
  XNOR2XL U588 ( .A(n31), .B(n220), .Y(SUM[9]) );
  XOR2XL U589 ( .A(n32), .B(n223), .Y(SUM[8]) );
  XNOR2XL U590 ( .A(n33), .B(n228), .Y(SUM[7]) );
  XOR2XL U591 ( .A(n34), .B(n231), .Y(SUM[6]) );
  XOR2XL U592 ( .A(n35), .B(n235), .Y(SUM[5]) );
  XNOR2XL U593 ( .A(n36), .B(n240), .Y(SUM[4]) );
  XOR2XL U594 ( .A(n37), .B(n243), .Y(SUM[3]) );
  XNOR2X1 U595 ( .A(n38), .B(n424), .Y(SUM[2]) );
  XNOR2X1 U596 ( .A(n39), .B(n254), .Y(SUM[1]) );
  NAND2BX1 U597 ( .AN(n255), .B(n256), .Y(n40) );
  NOR2X1 U598 ( .A(B[0]), .B(A[0]), .Y(n255) );
  INVX2 U599 ( .A(n40), .Y(SUM[0]) );
endmodule


module MMSA_DW01_add_43 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n63, n64, n65, n66, n67, n68, n69, n70, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n128, n129, n130, n131, n132, n133,
         n136, n137, n138, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n153, n155, n156, n157, n158, n160, n163,
         n164, n165, n166, n167, n169, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n201, n203, n204, n205, n206, n207, n209, n211, n212, n213,
         n214, n215, n217, n219, n220, n221, n222, n223, n225, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n237, n239, n240, n241,
         n242, n243, n245, n247, n253, n254, n255, n256, n270, n273, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435;

  AOI21X1 U27 ( .A0(n58), .A1(n86), .B0(n59), .Y(n57) );
  AOI21X1 U53 ( .A0(n86), .A1(n78), .B0(n79), .Y(n77) );
  AOI21X1 U116 ( .A0(n123), .A1(n143), .B0(n124), .Y(n122) );
  AOI21X1 U126 ( .A0(n143), .A1(n130), .B0(n131), .Y(n129) );
  AOI21X1 U138 ( .A0(n143), .A1(n270), .B0(n140), .Y(n138) );
  OAI21X2 U340 ( .A0(n109), .A1(n113), .B0(n110), .Y(n104) );
  NOR2X2 U341 ( .A(n80), .B(n73), .Y(n67) );
  NOR2X1 U342 ( .A(B[34]), .B(A[34]), .Y(n80) );
  NOR2X2 U343 ( .A(n60), .B(n53), .Y(n51) );
  AOI21XL U344 ( .A0(n104), .A1(n96), .B0(n97), .Y(n95) );
  NOR2X2 U345 ( .A(B[35]), .B(A[35]), .Y(n73) );
  OAI21X1 U346 ( .A0(n73), .A1(n81), .B0(n74), .Y(n68) );
  NAND2X1 U347 ( .A(B[34]), .B(A[34]), .Y(n81) );
  OAI21X4 U348 ( .A0(n151), .A1(n147), .B0(n148), .Y(n146) );
  AOI21X2 U349 ( .A0(n429), .A1(n160), .B0(n153), .Y(n151) );
  AOI21X2 U350 ( .A0(n172), .A1(n426), .B0(n169), .Y(n167) );
  OAI21X2 U351 ( .A0(n187), .A1(n185), .B0(n186), .Y(n184) );
  OAI21X2 U352 ( .A0(n165), .A1(n167), .B0(n166), .Y(n164) );
  NOR2X1 U353 ( .A(B[15]), .B(A[15]), .Y(n193) );
  NOR2X1 U354 ( .A(n112), .B(n109), .Y(n103) );
  OAI21X1 U355 ( .A0(n116), .A1(n144), .B0(n117), .Y(n115) );
  NOR2X1 U356 ( .A(B[10]), .B(A[10]), .Y(n213) );
  NOR2X1 U357 ( .A(B[12]), .B(A[12]), .Y(n205) );
  NOR2X1 U358 ( .A(B[20]), .B(A[20]), .Y(n173) );
  OAI21X2 U359 ( .A0(n173), .A1(n423), .B0(n174), .Y(n172) );
  AOI21X1 U360 ( .A0(n176), .A1(n184), .B0(n177), .Y(n423) );
  NOR2X1 U361 ( .A(B[28]), .B(A[28]), .Y(n125) );
  NOR2X1 U362 ( .A(B[30]), .B(A[30]), .Y(n112) );
  NOR2X1 U363 ( .A(B[17]), .B(A[17]), .Y(n185) );
  NOR2X1 U364 ( .A(B[25]), .B(A[25]), .Y(n147) );
  NOR2X1 U365 ( .A(B[33]), .B(A[33]), .Y(n91) );
  AOI21X1 U366 ( .A0(n89), .A1(n104), .B0(n90), .Y(n84) );
  AOI21XL U367 ( .A0(n86), .A1(n67), .B0(n68), .Y(n66) );
  AOI21XL U368 ( .A0(n51), .A1(n68), .B0(n52), .Y(n50) );
  AOI21X1 U369 ( .A0(n131), .A1(n118), .B0(n119), .Y(n117) );
  AOI21XL U370 ( .A0(n176), .A1(n184), .B0(n177), .Y(n175) );
  NAND2X1 U371 ( .A(n130), .B(n118), .Y(n116) );
  NOR2X1 U372 ( .A(n125), .B(n120), .Y(n118) );
  OR2XL U373 ( .A(B[11]), .B(A[11]), .Y(n431) );
  NAND2XL U374 ( .A(B[8]), .B(A[8]), .Y(n222) );
  OAI21XL U375 ( .A0(n114), .A1(n65), .B0(n66), .Y(n64) );
  OAI21XL U376 ( .A0(n114), .A1(n76), .B0(n77), .Y(n75) );
  CLKINVXL U377 ( .A(n81), .Y(n79) );
  NAND2XL U378 ( .A(n85), .B(n67), .Y(n65) );
  INVX1 U379 ( .A(n115), .Y(n114) );
  OAI21X1 U380 ( .A0(n91), .A1(n99), .B0(n92), .Y(n90) );
  OAI21X1 U381 ( .A0(n114), .A1(n56), .B0(n57), .Y(n55) );
  NOR2X1 U382 ( .A(n91), .B(n98), .Y(n89) );
  NOR2X1 U383 ( .A(B[19]), .B(A[19]), .Y(n178) );
  NOR2X1 U384 ( .A(B[27]), .B(A[27]), .Y(n136) );
  NAND2BX1 U385 ( .AN(n41), .B(n42), .Y(n1) );
  OR2X1 U386 ( .A(B[7]), .B(A[7]), .Y(n430) );
  OR2X1 U387 ( .A(B[9]), .B(A[9]), .Y(n433) );
  OAI21XL U388 ( .A0(n114), .A1(n101), .B0(n102), .Y(n100) );
  CLKINVX1 U389 ( .A(n232), .Y(n231) );
  NAND2BX1 U390 ( .AN(n120), .B(n121), .Y(n11) );
  OR2XL U391 ( .A(B[24]), .B(A[24]), .Y(n429) );
  NAND2X1 U392 ( .A(B[10]), .B(A[10]), .Y(n214) );
  NAND2X1 U393 ( .A(n89), .B(n103), .Y(n83) );
  CLKINVXL U394 ( .A(n84), .Y(n86) );
  CLKINVXL U395 ( .A(n104), .Y(n102) );
  CLKINVXL U396 ( .A(n144), .Y(n143) );
  CLKINVXL U397 ( .A(n164), .Y(n163) );
  OAI21XL U398 ( .A0(n163), .A1(n150), .B0(n151), .Y(n149) );
  NOR2X2 U399 ( .A(n141), .B(n136), .Y(n130) );
  CLKINVXL U400 ( .A(n99), .Y(n97) );
  CLKINVXL U401 ( .A(n98), .Y(n96) );
  NAND2XL U402 ( .A(n96), .B(n99), .Y(n8) );
  AOI21X1 U403 ( .A0(n188), .A1(n196), .B0(n189), .Y(n187) );
  OAI21XL U404 ( .A0(n53), .A1(n63), .B0(n54), .Y(n52) );
  OAI21XL U405 ( .A0(n70), .A1(n60), .B0(n63), .Y(n59) );
  CLKINVX2 U406 ( .A(n157), .Y(n273) );
  OAI21XL U407 ( .A0(n163), .A1(n157), .B0(n158), .Y(n156) );
  CLKINVXL U408 ( .A(n141), .Y(n270) );
  CLKINVXL U409 ( .A(n80), .Y(n78) );
  NAND2BXL U410 ( .AN(n173), .B(n174), .Y(n20) );
  NAND2BXL U411 ( .AN(n178), .B(n179), .Y(n21) );
  NAND2XL U412 ( .A(n273), .B(n158), .Y(n17) );
  NAND2BXL U413 ( .AN(n205), .B(n206), .Y(n28) );
  NAND2XL U414 ( .A(B[27]), .B(A[27]), .Y(n137) );
  NAND2XL U415 ( .A(B[26]), .B(A[26]), .Y(n142) );
  NAND2XL U416 ( .A(B[30]), .B(A[30]), .Y(n113) );
  NAND2XL U417 ( .A(B[28]), .B(A[28]), .Y(n128) );
  NAND2XL U418 ( .A(B[18]), .B(A[18]), .Y(n182) );
  NAND2XL U419 ( .A(B[15]), .B(A[15]), .Y(n194) );
  NOR2X1 U420 ( .A(B[29]), .B(A[29]), .Y(n120) );
  OR2XL U421 ( .A(B[13]), .B(A[13]), .Y(n425) );
  NAND2XL U422 ( .A(B[21]), .B(A[21]), .Y(n171) );
  NAND2XL U423 ( .A(B[13]), .B(A[13]), .Y(n203) );
  NAND2XL U424 ( .A(B[24]), .B(A[24]), .Y(n155) );
  OR2XL U425 ( .A(B[21]), .B(A[21]), .Y(n426) );
  NAND2XL U426 ( .A(B[17]), .B(A[17]), .Y(n186) );
  NAND2XL U427 ( .A(B[11]), .B(A[11]), .Y(n211) );
  NAND2XL U428 ( .A(B[14]), .B(A[14]), .Y(n198) );
  NAND2XL U429 ( .A(B[23]), .B(A[23]), .Y(n158) );
  NAND2XL U430 ( .A(B[22]), .B(A[22]), .Y(n166) );
  NAND2XL U431 ( .A(B[36]), .B(A[36]), .Y(n63) );
  NAND2XL U432 ( .A(B[7]), .B(A[7]), .Y(n227) );
  NAND2XL U433 ( .A(B[6]), .B(A[6]), .Y(n230) );
  NAND2XL U434 ( .A(B[9]), .B(A[9]), .Y(n219) );
  NAND2XL U435 ( .A(n434), .B(A[38]), .Y(n45) );
  NAND2XL U436 ( .A(B[5]), .B(A[5]), .Y(n234) );
  OR2XL U437 ( .A(B[4]), .B(A[4]), .Y(n428) );
  NAND2XL U438 ( .A(B[4]), .B(A[4]), .Y(n239) );
  NOR2X1 U439 ( .A(B[3]), .B(A[3]), .Y(n241) );
  NAND2XL U440 ( .A(B[3]), .B(A[3]), .Y(n242) );
  INVX2 U441 ( .A(n435), .Y(n434) );
  INVX2 U442 ( .A(B[38]), .Y(n435) );
  INVX2 U443 ( .A(n83), .Y(n85) );
  AOI21X1 U444 ( .A0(n115), .A1(n47), .B0(n48), .Y(n46) );
  NOR2X1 U445 ( .A(n49), .B(n83), .Y(n47) );
  OAI21X1 U446 ( .A0(n84), .A1(n49), .B0(n50), .Y(n48) );
  NAND2X1 U447 ( .A(n67), .B(n51), .Y(n49) );
  INVX2 U448 ( .A(n67), .Y(n69) );
  OAI21XL U449 ( .A0(n114), .A1(n83), .B0(n84), .Y(n82) );
  CLKINVXL U450 ( .A(n103), .Y(n101) );
  INVX2 U451 ( .A(n130), .Y(n132) );
  INVX2 U452 ( .A(n184), .Y(n183) );
  INVX2 U453 ( .A(n196), .Y(n195) );
  OAI21X1 U454 ( .A0(n46), .A1(n44), .B0(n45), .Y(n43) );
  NAND2XL U455 ( .A(n58), .B(n85), .Y(n56) );
  NOR2X1 U456 ( .A(n69), .B(n60), .Y(n58) );
  CLKINVXL U457 ( .A(n68), .Y(n70) );
  OAI21X1 U458 ( .A0(n178), .A1(n182), .B0(n179), .Y(n177) );
  INVX2 U459 ( .A(n171), .Y(n169) );
  AOI21X2 U460 ( .A0(n145), .A1(n164), .B0(n146), .Y(n144) );
  NOR2X1 U461 ( .A(n150), .B(n147), .Y(n145) );
  OAI21X1 U462 ( .A0(n199), .A1(n197), .B0(n198), .Y(n196) );
  OAI21X1 U463 ( .A0(n190), .A1(n194), .B0(n191), .Y(n189) );
  NOR2X1 U464 ( .A(n193), .B(n190), .Y(n188) );
  OAI21X1 U465 ( .A0(n205), .A1(n207), .B0(n206), .Y(n204) );
  AOI21X1 U466 ( .A0(n204), .A1(n425), .B0(n201), .Y(n199) );
  INVX2 U467 ( .A(n203), .Y(n201) );
  AOI21X1 U468 ( .A0(n428), .A1(n240), .B0(n237), .Y(n235) );
  INVX2 U469 ( .A(n239), .Y(n237) );
  AOI21X1 U470 ( .A0(n427), .A1(n424), .B0(n245), .Y(n243) );
  AOI21X1 U471 ( .A0(n220), .A1(n433), .B0(n217), .Y(n215) );
  INVX2 U472 ( .A(n219), .Y(n217) );
  AOI21X1 U473 ( .A0(n228), .A1(n430), .B0(n225), .Y(n223) );
  INVX2 U474 ( .A(n227), .Y(n225) );
  OAI21X1 U475 ( .A0(n221), .A1(n223), .B0(n222), .Y(n220) );
  OAI21X1 U476 ( .A0(n213), .A1(n215), .B0(n214), .Y(n212) );
  OAI21X1 U477 ( .A0(n229), .A1(n231), .B0(n230), .Y(n228) );
  OAI21X1 U478 ( .A0(n241), .A1(n243), .B0(n242), .Y(n240) );
  AOI21X1 U479 ( .A0(n431), .A1(n212), .B0(n209), .Y(n207) );
  INVX2 U480 ( .A(n211), .Y(n209) );
  OAI21X1 U481 ( .A0(n233), .A1(n235), .B0(n234), .Y(n232) );
  NAND2XL U482 ( .A(n85), .B(n78), .Y(n76) );
  OAI21X1 U483 ( .A0(n142), .A1(n136), .B0(n137), .Y(n131) );
  OAI21XL U484 ( .A0(n114), .A1(n112), .B0(n113), .Y(n111) );
  OAI21XL U485 ( .A0(n114), .A1(n94), .B0(n95), .Y(n93) );
  NAND2XL U486 ( .A(n103), .B(n96), .Y(n94) );
  INVX2 U487 ( .A(n155), .Y(n153) );
  INVX2 U488 ( .A(n158), .Y(n160) );
  OAI21XL U489 ( .A0(n133), .A1(n125), .B0(n128), .Y(n124) );
  NOR2X1 U490 ( .A(n132), .B(n125), .Y(n123) );
  CLKINVXL U491 ( .A(n131), .Y(n133) );
  INVX2 U492 ( .A(n142), .Y(n140) );
  OAI2BB1X1 U493 ( .A0N(n432), .A1N(n254), .B0(n253), .Y(n424) );
  OAI21X1 U494 ( .A0(n120), .A1(n128), .B0(n121), .Y(n119) );
  NAND2BX1 U495 ( .AN(n44), .B(n45), .Y(n2) );
  NAND2X1 U496 ( .A(n273), .B(n429), .Y(n150) );
  NAND2BX1 U497 ( .AN(n53), .B(n54), .Y(n3) );
  NAND2BX1 U498 ( .AN(n60), .B(n63), .Y(n4) );
  NAND2XL U499 ( .A(n78), .B(n81), .Y(n6) );
  NAND2BX1 U500 ( .AN(n73), .B(n74), .Y(n5) );
  NAND2BX1 U501 ( .AN(n91), .B(n92), .Y(n7) );
  NAND2BX1 U502 ( .AN(n125), .B(n128), .Y(n12) );
  INVX2 U503 ( .A(n256), .Y(n254) );
  NAND2BX1 U504 ( .AN(n112), .B(n113), .Y(n10) );
  NAND2BX1 U505 ( .AN(n147), .B(n148), .Y(n15) );
  NAND2BX1 U506 ( .AN(n109), .B(n110), .Y(n9) );
  NAND2X1 U507 ( .A(n270), .B(n142), .Y(n14) );
  NAND2BX1 U508 ( .AN(n136), .B(n137), .Y(n13) );
  NAND2X1 U509 ( .A(n426), .B(n171), .Y(n19) );
  NAND2X1 U510 ( .A(n429), .B(n155), .Y(n16) );
  NAND2BX1 U511 ( .AN(n165), .B(n166), .Y(n18) );
  NAND2BX1 U512 ( .AN(n181), .B(n182), .Y(n22) );
  NAND2BX1 U513 ( .AN(n185), .B(n186), .Y(n23) );
  OAI21XL U514 ( .A0(n195), .A1(n193), .B0(n194), .Y(n192) );
  NAND2BX1 U515 ( .AN(n197), .B(n198), .Y(n26) );
  NAND2BX1 U516 ( .AN(n190), .B(n191), .Y(n24) );
  NAND2BX1 U517 ( .AN(n193), .B(n194), .Y(n25) );
  NAND2X1 U518 ( .A(n425), .B(n203), .Y(n27) );
  NAND2X1 U519 ( .A(n431), .B(n211), .Y(n29) );
  NAND2BX1 U520 ( .AN(n213), .B(n214), .Y(n30) );
  NAND2X1 U521 ( .A(n433), .B(n219), .Y(n31) );
  NAND2BX1 U522 ( .AN(n221), .B(n222), .Y(n32) );
  NAND2X1 U523 ( .A(n430), .B(n227), .Y(n33) );
  NAND2BX1 U524 ( .AN(n229), .B(n230), .Y(n34) );
  NAND2BX1 U525 ( .AN(n233), .B(n234), .Y(n35) );
  NAND2X1 U526 ( .A(n428), .B(n239), .Y(n36) );
  NAND2BX1 U527 ( .AN(n241), .B(n242), .Y(n37) );
  NAND2XL U528 ( .A(n427), .B(n247), .Y(n38) );
  NAND2X1 U529 ( .A(n432), .B(n253), .Y(n39) );
  NOR2X1 U530 ( .A(B[37]), .B(A[37]), .Y(n53) );
  XNOR2X1 U531 ( .A(n43), .B(n1), .Y(SUM[39]) );
  NOR2X1 U532 ( .A(B[36]), .B(A[36]), .Y(n60) );
  XNOR2X1 U533 ( .A(n55), .B(n3), .Y(SUM[37]) );
  XOR2X1 U534 ( .A(n46), .B(n2), .Y(SUM[38]) );
  NOR2X1 U535 ( .A(B[31]), .B(A[31]), .Y(n109) );
  NAND2XL U536 ( .A(B[35]), .B(A[35]), .Y(n74) );
  NAND2XL U537 ( .A(B[37]), .B(A[37]), .Y(n54) );
  NOR2X1 U538 ( .A(B[18]), .B(A[18]), .Y(n181) );
  XNOR2X1 U539 ( .A(n82), .B(n6), .Y(SUM[34]) );
  NOR2X1 U540 ( .A(B[14]), .B(A[14]), .Y(n197) );
  NOR2X1 U541 ( .A(B[16]), .B(A[16]), .Y(n190) );
  XNOR2X1 U542 ( .A(n64), .B(n4), .Y(SUM[36]) );
  XNOR2X1 U543 ( .A(n75), .B(n5), .Y(SUM[35]) );
  XNOR2X1 U544 ( .A(n111), .B(n9), .Y(SUM[31]) );
  XNOR2X1 U545 ( .A(n100), .B(n8), .Y(SUM[32]) );
  XNOR2X1 U546 ( .A(n93), .B(n7), .Y(SUM[33]) );
  OR2X1 U547 ( .A(B[2]), .B(A[2]), .Y(n427) );
  NOR2X1 U548 ( .A(B[26]), .B(A[26]), .Y(n141) );
  XOR2X1 U549 ( .A(n122), .B(n11), .Y(SUM[29]) );
  NOR2X1 U550 ( .A(B[5]), .B(A[5]), .Y(n233) );
  XOR2X1 U551 ( .A(n129), .B(n12), .Y(SUM[28]) );
  XOR2X1 U552 ( .A(n138), .B(n13), .Y(SUM[27]) );
  XOR2X1 U553 ( .A(n114), .B(n10), .Y(SUM[30]) );
  NOR2X1 U554 ( .A(B[32]), .B(A[32]), .Y(n98) );
  OR2X1 U555 ( .A(B[1]), .B(A[1]), .Y(n432) );
  NOR2X1 U556 ( .A(B[6]), .B(A[6]), .Y(n229) );
  NOR2X1 U557 ( .A(n434), .B(A[38]), .Y(n44) );
  NAND2XL U558 ( .A(B[19]), .B(A[19]), .Y(n179) );
  NAND2X1 U559 ( .A(B[32]), .B(A[32]), .Y(n99) );
  NAND2XL U560 ( .A(B[12]), .B(A[12]), .Y(n206) );
  NAND2XL U561 ( .A(B[20]), .B(A[20]), .Y(n174) );
  NOR2X1 U562 ( .A(B[8]), .B(A[8]), .Y(n221) );
  NAND2XL U563 ( .A(B[29]), .B(A[29]), .Y(n121) );
  NAND2XL U564 ( .A(B[31]), .B(A[31]), .Y(n110) );
  NAND2XL U565 ( .A(n434), .B(A[39]), .Y(n42) );
  NOR2X1 U566 ( .A(n434), .B(A[39]), .Y(n41) );
  NAND2X1 U567 ( .A(B[1]), .B(A[1]), .Y(n253) );
  NAND2XL U568 ( .A(B[33]), .B(A[33]), .Y(n92) );
  NAND2XL U569 ( .A(B[16]), .B(A[16]), .Y(n191) );
  NOR2X1 U570 ( .A(B[23]), .B(A[23]), .Y(n157) );
  NAND2XL U571 ( .A(B[25]), .B(A[25]), .Y(n148) );
  XNOR2X1 U572 ( .A(n156), .B(n16), .Y(SUM[24]) );
  XNOR2X1 U573 ( .A(n149), .B(n15), .Y(SUM[25]) );
  XNOR2X1 U574 ( .A(n143), .B(n14), .Y(SUM[26]) );
  XOR2X1 U575 ( .A(n163), .B(n17), .Y(SUM[23]) );
  NOR2X1 U576 ( .A(B[22]), .B(A[22]), .Y(n165) );
  NAND2X1 U577 ( .A(B[0]), .B(A[0]), .Y(n256) );
  XOR2XL U578 ( .A(n18), .B(n167), .Y(SUM[22]) );
  XNOR2X1 U579 ( .A(n180), .B(n21), .Y(SUM[19]) );
  XNOR2X1 U580 ( .A(n172), .B(n19), .Y(SUM[21]) );
  XOR2XL U581 ( .A(n20), .B(n175), .Y(SUM[20]) );
  XOR2X1 U582 ( .A(n183), .B(n22), .Y(SUM[18]) );
  XOR2X1 U583 ( .A(n187), .B(n23), .Y(SUM[17]) );
  XNOR2X1 U584 ( .A(n192), .B(n24), .Y(SUM[16]) );
  XOR2X1 U585 ( .A(n25), .B(n195), .Y(SUM[15]) );
  XOR2XL U586 ( .A(n26), .B(n199), .Y(SUM[14]) );
  XNOR2XL U587 ( .A(n27), .B(n204), .Y(SUM[13]) );
  XOR2XL U588 ( .A(n28), .B(n207), .Y(SUM[12]) );
  XNOR2XL U589 ( .A(n29), .B(n212), .Y(SUM[11]) );
  XOR2XL U590 ( .A(n30), .B(n215), .Y(SUM[10]) );
  XNOR2XL U591 ( .A(n31), .B(n220), .Y(SUM[9]) );
  XOR2XL U592 ( .A(n32), .B(n223), .Y(SUM[8]) );
  XNOR2XL U593 ( .A(n33), .B(n228), .Y(SUM[7]) );
  XOR2XL U594 ( .A(n34), .B(n231), .Y(SUM[6]) );
  XOR2XL U595 ( .A(n35), .B(n235), .Y(SUM[5]) );
  XNOR2XL U596 ( .A(n36), .B(n240), .Y(SUM[4]) );
  XOR2XL U597 ( .A(n37), .B(n243), .Y(SUM[3]) );
  XNOR2XL U598 ( .A(n38), .B(n424), .Y(SUM[2]) );
  XNOR2X1 U599 ( .A(n39), .B(n254), .Y(SUM[1]) );
  NAND2BX1 U600 ( .AN(n255), .B(n256), .Y(n40) );
  NOR2X1 U601 ( .A(B[0]), .B(A[0]), .Y(n255) );
  INVX2 U602 ( .A(n40), .Y(SUM[0]) );
  NOR2X1 U603 ( .A(n181), .B(n178), .Y(n176) );
  OAI21XL U604 ( .A0(n183), .A1(n181), .B0(n182), .Y(n180) );
  INVX2 U605 ( .A(n247), .Y(n245) );
  NAND2XL U606 ( .A(B[2]), .B(A[2]), .Y(n247) );
endmodule


module MMSA_DW01_add_42 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n63, n64, n65, n66, n67, n68, n69, n70, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n128, n129, n130, n131, n133, n136,
         n137, n138, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n153, n155, n156, n157, n158, n160, n163, n164,
         n165, n166, n167, n169, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n201, n203, n204, n205, n206, n207, n209, n211, n212, n213, n214,
         n215, n217, n219, n220, n221, n222, n223, n225, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n237, n239, n240, n241, n242,
         n243, n245, n247, n253, n254, n255, n256, n270, n273, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436;

  AOI21X1 U17 ( .A0(n51), .A1(n68), .B0(n52), .Y(n50) );
  AOI21X1 U27 ( .A0(n58), .A1(n86), .B0(n59), .Y(n57) );
  NOR2X2 U34 ( .A(B[36]), .B(A[36]), .Y(n60) );
  AOI21X1 U39 ( .A0(n86), .A1(n67), .B0(n423), .Y(n66) );
  NOR2X2 U44 ( .A(n80), .B(n73), .Y(n67) );
  AOI21X1 U53 ( .A0(n86), .A1(n78), .B0(n79), .Y(n77) );
  AOI21X1 U77 ( .A0(n104), .A1(n96), .B0(n97), .Y(n95) );
  AOI21X1 U108 ( .A0(n131), .A1(n118), .B0(n119), .Y(n117) );
  AOI21X1 U116 ( .A0(n123), .A1(n143), .B0(n124), .Y(n122) );
  AOI21X1 U126 ( .A0(n143), .A1(n130), .B0(n131), .Y(n129) );
  AOI21X1 U138 ( .A0(n143), .A1(n270), .B0(n140), .Y(n138) );
  AOI21X1 U157 ( .A0(n426), .A1(n160), .B0(n153), .Y(n151) );
  AOI21X1 U196 ( .A0(n176), .A1(n184), .B0(n177), .Y(n175) );
  AOI21X1 U301 ( .A0(n429), .A1(n240), .B0(n237), .Y(n235) );
  OAI21X4 U340 ( .A0(n109), .A1(n113), .B0(n110), .Y(n104) );
  INVX1 U341 ( .A(n81), .Y(n79) );
  NOR2XL U342 ( .A(B[34]), .B(A[34]), .Y(n80) );
  OAI21X2 U343 ( .A0(n173), .A1(n175), .B0(n174), .Y(n172) );
  NOR2X1 U344 ( .A(n91), .B(n98), .Y(n89) );
  NOR2X1 U345 ( .A(n112), .B(n109), .Y(n103) );
  NOR2X1 U346 ( .A(n60), .B(n53), .Y(n51) );
  AOI21X1 U347 ( .A0(n89), .A1(n104), .B0(n90), .Y(n84) );
  OAI21X1 U348 ( .A0(n116), .A1(n424), .B0(n117), .Y(n115) );
  AOI21XL U349 ( .A0(n145), .A1(n164), .B0(n146), .Y(n424) );
  NOR2X1 U350 ( .A(n125), .B(n120), .Y(n118) );
  NAND2X1 U351 ( .A(B[23]), .B(A[23]), .Y(n158) );
  NOR2X1 U352 ( .A(B[28]), .B(A[28]), .Y(n125) );
  NOR2X1 U353 ( .A(B[30]), .B(A[30]), .Y(n112) );
  NOR2X1 U354 ( .A(B[29]), .B(A[29]), .Y(n120) );
  NOR2X1 U355 ( .A(B[33]), .B(A[33]), .Y(n91) );
  NAND2X1 U356 ( .A(n67), .B(n51), .Y(n49) );
  OAI21X2 U357 ( .A0(n165), .A1(n167), .B0(n166), .Y(n164) );
  CLKINVXL U358 ( .A(n70), .Y(n423) );
  AOI21XL U359 ( .A0(n145), .A1(n164), .B0(n146), .Y(n144) );
  OAI21X1 U360 ( .A0(n151), .A1(n147), .B0(n148), .Y(n146) );
  OR2X1 U361 ( .A(B[24]), .B(A[24]), .Y(n426) );
  NAND2BX1 U362 ( .AN(n41), .B(n42), .Y(n1) );
  OAI21XL U363 ( .A0(n114), .A1(n101), .B0(n102), .Y(n100) );
  OAI21XL U364 ( .A0(n114), .A1(n56), .B0(n57), .Y(n55) );
  NOR2X1 U365 ( .A(B[35]), .B(A[35]), .Y(n73) );
  OR2X1 U366 ( .A(B[4]), .B(A[4]), .Y(n429) );
  CLKINVXL U367 ( .A(n83), .Y(n85) );
  CLKINVXL U368 ( .A(n84), .Y(n86) );
  INVX1 U369 ( .A(n115), .Y(n114) );
  CLKINVXL U370 ( .A(n131), .Y(n133) );
  CLKINVXL U371 ( .A(n184), .Y(n183) );
  CLKINVXL U372 ( .A(n196), .Y(n195) );
  CLKINVXL U373 ( .A(n99), .Y(n97) );
  CLKINVXL U374 ( .A(n98), .Y(n96) );
  NAND2XL U375 ( .A(n96), .B(n99), .Y(n8) );
  OAI21X1 U376 ( .A0(n120), .A1(n128), .B0(n121), .Y(n119) );
  NOR2BXL U377 ( .AN(n130), .B(n125), .Y(n123) );
  OAI21XL U378 ( .A0(n53), .A1(n63), .B0(n54), .Y(n52) );
  CLKINVX1 U379 ( .A(n227), .Y(n225) );
  CLKINVX2 U380 ( .A(n157), .Y(n273) );
  CLKINVXL U381 ( .A(n141), .Y(n270) );
  NAND2BXL U382 ( .AN(n73), .B(n74), .Y(n5) );
  INVX1 U383 ( .A(n232), .Y(n231) );
  NAND2BXL U384 ( .AN(n125), .B(n128), .Y(n12) );
  NAND2BXL U385 ( .AN(n112), .B(n113), .Y(n10) );
  NAND2XL U386 ( .A(n273), .B(n158), .Y(n17) );
  OAI21XL U387 ( .A0(n183), .A1(n181), .B0(n182), .Y(n180) );
  OAI21XL U388 ( .A0(n195), .A1(n193), .B0(n194), .Y(n192) );
  NAND2XL U389 ( .A(n430), .B(n211), .Y(n29) );
  NAND2XL U390 ( .A(n433), .B(n219), .Y(n31) );
  NAND2XL U391 ( .A(n432), .B(n227), .Y(n33) );
  NAND2XL U392 ( .A(B[26]), .B(A[26]), .Y(n142) );
  NAND2XL U393 ( .A(B[18]), .B(A[18]), .Y(n182) );
  NAND2XL U394 ( .A(B[15]), .B(A[15]), .Y(n194) );
  OR2XL U395 ( .A(B[13]), .B(A[13]), .Y(n427) );
  NAND2XL U396 ( .A(B[13]), .B(A[13]), .Y(n203) );
  OR2XL U397 ( .A(B[21]), .B(A[21]), .Y(n428) );
  NAND2XL U398 ( .A(B[34]), .B(A[34]), .Y(n81) );
  NAND2XL U399 ( .A(B[21]), .B(A[21]), .Y(n171) );
  NAND2XL U400 ( .A(B[36]), .B(A[36]), .Y(n63) );
  NAND2XL U401 ( .A(B[24]), .B(A[24]), .Y(n155) );
  OR2XL U402 ( .A(B[7]), .B(A[7]), .Y(n432) );
  NAND2XL U403 ( .A(B[22]), .B(A[22]), .Y(n166) );
  OR2XL U404 ( .A(B[9]), .B(A[9]), .Y(n433) );
  NAND2XL U405 ( .A(n435), .B(A[38]), .Y(n45) );
  NAND2XL U406 ( .A(B[4]), .B(A[4]), .Y(n239) );
  NAND2XL U407 ( .A(B[3]), .B(A[3]), .Y(n242) );
  INVX2 U408 ( .A(n436), .Y(n435) );
  INVX2 U409 ( .A(B[38]), .Y(n436) );
  AOI21X1 U410 ( .A0(n115), .A1(n47), .B0(n48), .Y(n46) );
  OAI21X1 U411 ( .A0(n84), .A1(n49), .B0(n50), .Y(n48) );
  NOR2X1 U412 ( .A(n49), .B(n83), .Y(n47) );
  CLKINVXL U413 ( .A(n67), .Y(n69) );
  OAI21X1 U414 ( .A0(n114), .A1(n65), .B0(n66), .Y(n64) );
  NAND2XL U415 ( .A(n85), .B(n67), .Y(n65) );
  NAND2X1 U416 ( .A(n89), .B(n103), .Y(n83) );
  OAI21XL U417 ( .A0(n114), .A1(n83), .B0(n84), .Y(n82) );
  INVX2 U418 ( .A(n104), .Y(n102) );
  CLKINVXL U419 ( .A(n103), .Y(n101) );
  INVX2 U420 ( .A(n144), .Y(n143) );
  INVX2 U421 ( .A(n164), .Y(n163) );
  OAI21X1 U422 ( .A0(n163), .A1(n150), .B0(n151), .Y(n149) );
  OAI21X1 U423 ( .A0(n46), .A1(n44), .B0(n45), .Y(n43) );
  NAND2XL U424 ( .A(n58), .B(n85), .Y(n56) );
  NOR2X1 U425 ( .A(n69), .B(n60), .Y(n58) );
  OAI21X1 U426 ( .A0(n73), .A1(n81), .B0(n74), .Y(n68) );
  OAI21XL U427 ( .A0(n70), .A1(n60), .B0(n63), .Y(n59) );
  CLKINVXL U428 ( .A(n68), .Y(n70) );
  OAI21X1 U429 ( .A0(n91), .A1(n99), .B0(n92), .Y(n90) );
  NAND2X1 U430 ( .A(n130), .B(n118), .Y(n116) );
  OAI21XL U431 ( .A0(n114), .A1(n76), .B0(n77), .Y(n75) );
  NAND2XL U432 ( .A(n85), .B(n78), .Y(n76) );
  OAI21X1 U433 ( .A0(n178), .A1(n182), .B0(n179), .Y(n177) );
  NOR2X1 U434 ( .A(n181), .B(n178), .Y(n176) );
  NOR2X1 U435 ( .A(n150), .B(n147), .Y(n145) );
  AOI21X1 U436 ( .A0(n188), .A1(n196), .B0(n189), .Y(n187) );
  OAI21X1 U437 ( .A0(n190), .A1(n194), .B0(n191), .Y(n189) );
  NOR2X1 U438 ( .A(n193), .B(n190), .Y(n188) );
  OAI21X1 U439 ( .A0(n187), .A1(n185), .B0(n186), .Y(n184) );
  AOI21X1 U440 ( .A0(n172), .A1(n428), .B0(n169), .Y(n167) );
  INVX2 U441 ( .A(n171), .Y(n169) );
  OAI21XL U442 ( .A0(n114), .A1(n112), .B0(n113), .Y(n111) );
  OAI21XL U443 ( .A0(n114), .A1(n94), .B0(n95), .Y(n93) );
  NAND2XL U444 ( .A(n103), .B(n96), .Y(n94) );
  OAI21X1 U445 ( .A0(n199), .A1(n197), .B0(n198), .Y(n196) );
  OAI21X1 U446 ( .A0(n142), .A1(n136), .B0(n137), .Y(n131) );
  OAI21XL U447 ( .A0(n133), .A1(n125), .B0(n128), .Y(n124) );
  INVX2 U448 ( .A(n142), .Y(n140) );
  AOI21X1 U449 ( .A0(n204), .A1(n427), .B0(n201), .Y(n199) );
  INVX2 U450 ( .A(n203), .Y(n201) );
  AOI21X1 U451 ( .A0(n430), .A1(n212), .B0(n209), .Y(n207) );
  INVX2 U452 ( .A(n211), .Y(n209) );
  AOI21X1 U453 ( .A0(n228), .A1(n432), .B0(n225), .Y(n223) );
  OAI21X1 U454 ( .A0(n221), .A1(n223), .B0(n222), .Y(n220) );
  OAI21X1 U455 ( .A0(n205), .A1(n207), .B0(n206), .Y(n204) );
  INVX2 U456 ( .A(n239), .Y(n237) );
  OAI21X1 U457 ( .A0(n229), .A1(n231), .B0(n230), .Y(n228) );
  OAI21X1 U458 ( .A0(n213), .A1(n215), .B0(n214), .Y(n212) );
  OAI21X1 U459 ( .A0(n241), .A1(n243), .B0(n242), .Y(n240) );
  AOI21X1 U460 ( .A0(n431), .A1(n425), .B0(n245), .Y(n243) );
  INVX2 U461 ( .A(n247), .Y(n245) );
  AOI21X1 U462 ( .A0(n220), .A1(n433), .B0(n217), .Y(n215) );
  INVX2 U463 ( .A(n219), .Y(n217) );
  OAI21X1 U464 ( .A0(n233), .A1(n235), .B0(n234), .Y(n232) );
  NOR2X1 U465 ( .A(n141), .B(n136), .Y(n130) );
  INVX2 U466 ( .A(n155), .Y(n153) );
  INVX2 U467 ( .A(n158), .Y(n160) );
  CLKINVXL U468 ( .A(n80), .Y(n78) );
  NAND2BX1 U469 ( .AN(n44), .B(n45), .Y(n2) );
  NAND2BX1 U470 ( .AN(n53), .B(n54), .Y(n3) );
  NAND2BX1 U471 ( .AN(n60), .B(n63), .Y(n4) );
  NAND2X1 U472 ( .A(n273), .B(n426), .Y(n150) );
  NAND2XL U473 ( .A(n78), .B(n81), .Y(n6) );
  OAI2BB1X1 U474 ( .A0N(n434), .A1N(n254), .B0(n253), .Y(n425) );
  OAI21X1 U475 ( .A0(n163), .A1(n157), .B0(n158), .Y(n156) );
  NAND2BX1 U476 ( .AN(n136), .B(n137), .Y(n13) );
  NAND2BX1 U477 ( .AN(n120), .B(n121), .Y(n11) );
  NAND2BX1 U478 ( .AN(n91), .B(n92), .Y(n7) );
  NAND2X1 U479 ( .A(n270), .B(n142), .Y(n14) );
  NAND2BX1 U480 ( .AN(n109), .B(n110), .Y(n9) );
  NAND2BX1 U481 ( .AN(n147), .B(n148), .Y(n15) );
  INVX2 U482 ( .A(n256), .Y(n254) );
  NAND2X1 U483 ( .A(n428), .B(n171), .Y(n19) );
  NAND2BX1 U484 ( .AN(n173), .B(n174), .Y(n20) );
  NAND2BX1 U485 ( .AN(n165), .B(n166), .Y(n18) );
  NAND2X1 U486 ( .A(n426), .B(n155), .Y(n16) );
  NAND2BX1 U487 ( .AN(n181), .B(n182), .Y(n22) );
  NAND2BX1 U488 ( .AN(n178), .B(n179), .Y(n21) );
  NAND2BX1 U489 ( .AN(n185), .B(n186), .Y(n23) );
  NAND2BX1 U490 ( .AN(n197), .B(n198), .Y(n26) );
  NAND2BX1 U491 ( .AN(n190), .B(n191), .Y(n24) );
  NAND2BX1 U492 ( .AN(n193), .B(n194), .Y(n25) );
  NAND2X1 U493 ( .A(n427), .B(n203), .Y(n27) );
  NAND2BX1 U494 ( .AN(n205), .B(n206), .Y(n28) );
  NAND2BX1 U495 ( .AN(n213), .B(n214), .Y(n30) );
  NAND2BX1 U496 ( .AN(n221), .B(n222), .Y(n32) );
  NAND2BX1 U497 ( .AN(n229), .B(n230), .Y(n34) );
  NAND2BX1 U498 ( .AN(n233), .B(n234), .Y(n35) );
  NAND2X1 U499 ( .A(n429), .B(n239), .Y(n36) );
  NAND2BX1 U500 ( .AN(n241), .B(n242), .Y(n37) );
  NAND2XL U501 ( .A(n431), .B(n247), .Y(n38) );
  NAND2X1 U502 ( .A(n434), .B(n253), .Y(n39) );
  XNOR2X1 U503 ( .A(n43), .B(n1), .Y(SUM[39]) );
  XNOR2X1 U504 ( .A(n55), .B(n3), .Y(SUM[37]) );
  NOR2X1 U505 ( .A(B[37]), .B(A[37]), .Y(n53) );
  XOR2X1 U506 ( .A(n46), .B(n2), .Y(SUM[38]) );
  XNOR2X1 U507 ( .A(n64), .B(n4), .Y(SUM[36]) );
  NOR2X1 U508 ( .A(B[31]), .B(A[31]), .Y(n109) );
  NAND2XL U509 ( .A(B[35]), .B(A[35]), .Y(n74) );
  XNOR2X1 U510 ( .A(n75), .B(n5), .Y(SUM[35]) );
  NAND2XL U511 ( .A(B[37]), .B(A[37]), .Y(n54) );
  XNOR2X1 U512 ( .A(n100), .B(n8), .Y(SUM[32]) );
  NOR2X1 U513 ( .A(B[16]), .B(A[16]), .Y(n190) );
  XNOR2X1 U514 ( .A(n111), .B(n9), .Y(SUM[31]) );
  XNOR2X1 U515 ( .A(n93), .B(n7), .Y(SUM[33]) );
  XNOR2X1 U516 ( .A(n82), .B(n6), .Y(SUM[34]) );
  NOR2X1 U517 ( .A(B[14]), .B(A[14]), .Y(n197) );
  NOR2X1 U518 ( .A(B[19]), .B(A[19]), .Y(n178) );
  NOR2X1 U519 ( .A(B[20]), .B(A[20]), .Y(n173) );
  NOR2X1 U520 ( .A(B[18]), .B(A[18]), .Y(n181) );
  NOR2X1 U521 ( .A(B[27]), .B(A[27]), .Y(n136) );
  XOR2X1 U522 ( .A(n122), .B(n11), .Y(SUM[29]) );
  XOR2X1 U523 ( .A(n114), .B(n10), .Y(SUM[30]) );
  NOR2X1 U524 ( .A(B[15]), .B(A[15]), .Y(n193) );
  XOR2X1 U525 ( .A(n129), .B(n12), .Y(SUM[28]) );
  XOR2X1 U526 ( .A(n138), .B(n13), .Y(SUM[27]) );
  NOR2X1 U527 ( .A(B[32]), .B(A[32]), .Y(n98) );
  NOR2X1 U528 ( .A(B[12]), .B(A[12]), .Y(n205) );
  NOR2X1 U529 ( .A(B[26]), .B(A[26]), .Y(n141) );
  NOR2X1 U530 ( .A(B[17]), .B(A[17]), .Y(n185) );
  NAND2XL U531 ( .A(B[14]), .B(A[14]), .Y(n198) );
  NAND2XL U532 ( .A(B[20]), .B(A[20]), .Y(n174) );
  NAND2XL U533 ( .A(B[19]), .B(A[19]), .Y(n179) );
  NAND2XL U534 ( .A(B[27]), .B(A[27]), .Y(n137) );
  NOR2X1 U535 ( .A(B[5]), .B(A[5]), .Y(n233) );
  NAND2XL U536 ( .A(B[28]), .B(A[28]), .Y(n128) );
  NAND2X1 U537 ( .A(B[30]), .B(A[30]), .Y(n113) );
  NOR2X1 U538 ( .A(n435), .B(A[38]), .Y(n44) );
  NOR2X1 U539 ( .A(B[25]), .B(A[25]), .Y(n147) );
  OR2XL U540 ( .A(B[11]), .B(A[11]), .Y(n430) );
  NAND2XL U541 ( .A(B[16]), .B(A[16]), .Y(n191) );
  NOR2X1 U542 ( .A(B[6]), .B(A[6]), .Y(n229) );
  NAND2XL U543 ( .A(B[12]), .B(A[12]), .Y(n206) );
  NAND2X1 U544 ( .A(B[32]), .B(A[32]), .Y(n99) );
  NOR2X1 U545 ( .A(B[10]), .B(A[10]), .Y(n213) );
  NAND2XL U546 ( .A(B[29]), .B(A[29]), .Y(n121) );
  NAND2X1 U547 ( .A(n435), .B(A[39]), .Y(n42) );
  NOR2X1 U548 ( .A(n435), .B(A[39]), .Y(n41) );
  OR2XL U549 ( .A(B[2]), .B(A[2]), .Y(n431) );
  NAND2XL U550 ( .A(B[33]), .B(A[33]), .Y(n92) );
  NAND2XL U551 ( .A(B[31]), .B(A[31]), .Y(n110) );
  NAND2XL U552 ( .A(B[17]), .B(A[17]), .Y(n186) );
  NAND2XL U553 ( .A(B[11]), .B(A[11]), .Y(n211) );
  NAND2XL U554 ( .A(B[25]), .B(A[25]), .Y(n148) );
  NAND2XL U555 ( .A(B[5]), .B(A[5]), .Y(n234) );
  NOR2X1 U556 ( .A(B[23]), .B(A[23]), .Y(n157) );
  NOR2X1 U557 ( .A(B[3]), .B(A[3]), .Y(n241) );
  NAND2XL U558 ( .A(B[7]), .B(A[7]), .Y(n227) );
  NAND2XL U559 ( .A(B[6]), .B(A[6]), .Y(n230) );
  NAND2XL U560 ( .A(B[10]), .B(A[10]), .Y(n214) );
  XNOR2X1 U561 ( .A(n143), .B(n14), .Y(SUM[26]) );
  NOR2X1 U562 ( .A(B[8]), .B(A[8]), .Y(n221) );
  OR2XL U563 ( .A(B[1]), .B(A[1]), .Y(n434) );
  NAND2XL U564 ( .A(B[9]), .B(A[9]), .Y(n219) );
  XNOR2X1 U565 ( .A(n156), .B(n16), .Y(SUM[24]) );
  XNOR2X1 U566 ( .A(n149), .B(n15), .Y(SUM[25]) );
  NOR2X1 U567 ( .A(B[22]), .B(A[22]), .Y(n165) );
  NAND2XL U568 ( .A(B[1]), .B(A[1]), .Y(n253) );
  NAND2XL U569 ( .A(B[8]), .B(A[8]), .Y(n222) );
  XOR2X1 U570 ( .A(n163), .B(n17), .Y(SUM[23]) );
  NAND2X1 U571 ( .A(B[0]), .B(A[0]), .Y(n256) );
  XNOR2X1 U572 ( .A(n180), .B(n21), .Y(SUM[19]) );
  XOR2X1 U573 ( .A(n183), .B(n22), .Y(SUM[18]) );
  XOR2X1 U574 ( .A(n187), .B(n23), .Y(SUM[17]) );
  XNOR2X1 U575 ( .A(n192), .B(n24), .Y(SUM[16]) );
  XOR2X1 U576 ( .A(n25), .B(n195), .Y(SUM[15]) );
  XOR2XL U577 ( .A(n26), .B(n199), .Y(SUM[14]) );
  XNOR2XL U578 ( .A(n27), .B(n204), .Y(SUM[13]) );
  XOR2XL U579 ( .A(n28), .B(n207), .Y(SUM[12]) );
  XNOR2XL U580 ( .A(n29), .B(n212), .Y(SUM[11]) );
  XNOR2XL U581 ( .A(n31), .B(n220), .Y(SUM[9]) );
  XOR2XL U582 ( .A(n32), .B(n223), .Y(SUM[8]) );
  XNOR2XL U583 ( .A(n33), .B(n228), .Y(SUM[7]) );
  XOR2XL U584 ( .A(n34), .B(n231), .Y(SUM[6]) );
  XNOR2XL U585 ( .A(n36), .B(n240), .Y(SUM[4]) );
  XNOR2X1 U586 ( .A(n38), .B(n425), .Y(SUM[2]) );
  XNOR2X1 U587 ( .A(n39), .B(n254), .Y(SUM[1]) );
  NAND2BX1 U588 ( .AN(n255), .B(n256), .Y(n40) );
  NOR2X1 U589 ( .A(B[0]), .B(A[0]), .Y(n255) );
  INVX2 U590 ( .A(n40), .Y(SUM[0]) );
  XOR2XL U591 ( .A(n18), .B(n167), .Y(SUM[22]) );
  XNOR2X1 U592 ( .A(n172), .B(n19), .Y(SUM[21]) );
  XOR2XL U593 ( .A(n20), .B(n175), .Y(SUM[20]) );
  XOR2XL U594 ( .A(n30), .B(n215), .Y(SUM[10]) );
  XOR2XL U595 ( .A(n35), .B(n235), .Y(SUM[5]) );
  XOR2XL U596 ( .A(n37), .B(n243), .Y(SUM[3]) );
  NAND2XL U597 ( .A(B[2]), .B(A[2]), .Y(n247) );
endmodule


module MMSA_DW01_add_41 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n63, n64, n65, n66, n67, n68, n69, n70, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n128, n129, n130, n131, n132, n133,
         n136, n137, n138, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n153, n155, n156, n157, n158, n160, n163,
         n164, n165, n166, n167, n169, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n201, n203, n204, n205, n206, n207, n209, n211, n212, n213,
         n214, n215, n217, n219, n220, n221, n222, n223, n225, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n237, n239, n240, n241,
         n242, n243, n245, n247, n253, n254, n255, n256, n270, n273, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438;

  AOI21X1 U27 ( .A0(n58), .A1(n86), .B0(n59), .Y(n57) );
  AOI21X1 U53 ( .A0(n86), .A1(n78), .B0(n79), .Y(n77) );
  AOI21X1 U77 ( .A0(n104), .A1(n96), .B0(n97), .Y(n95) );
  AOI21X1 U126 ( .A0(n143), .A1(n130), .B0(n131), .Y(n129) );
  NOR2X2 U135 ( .A(B[27]), .B(A[27]), .Y(n136) );
  AOI21X1 U157 ( .A0(n429), .A1(n160), .B0(n153), .Y(n151) );
  AOI21X1 U238 ( .A0(n204), .A1(n430), .B0(n201), .Y(n199) );
  AOI21X1 U252 ( .A0(n433), .A1(n212), .B0(n209), .Y(n207) );
  AOI21X1 U315 ( .A0(n434), .A1(n427), .B0(n245), .Y(n243) );
  NOR2XL U340 ( .A(B[34]), .B(A[34]), .Y(n80) );
  NOR2X2 U341 ( .A(B[37]), .B(A[37]), .Y(n53) );
  NOR2X2 U342 ( .A(B[36]), .B(A[36]), .Y(n60) );
  NOR2X2 U343 ( .A(B[33]), .B(A[33]), .Y(n91) );
  NOR2X2 U344 ( .A(B[31]), .B(A[31]), .Y(n109) );
  NAND2X1 U345 ( .A(n423), .B(n424), .Y(n425) );
  NAND2X1 U346 ( .A(n425), .B(n50), .Y(n48) );
  CLKINVXL U347 ( .A(n84), .Y(n423) );
  CLKINVX2 U348 ( .A(n49), .Y(n424) );
  AOI21XL U349 ( .A0(n51), .A1(n68), .B0(n52), .Y(n50) );
  INVX1 U350 ( .A(n67), .Y(n69) );
  NOR2X2 U351 ( .A(n80), .B(n73), .Y(n67) );
  OAI21X1 U352 ( .A0(n165), .A1(n167), .B0(n166), .Y(n164) );
  OAI21X1 U353 ( .A0(n151), .A1(n147), .B0(n148), .Y(n146) );
  NOR2X1 U354 ( .A(n91), .B(n98), .Y(n89) );
  NOR2X1 U355 ( .A(B[18]), .B(A[18]), .Y(n181) );
  NOR2X1 U356 ( .A(B[19]), .B(A[19]), .Y(n178) );
  NOR2X1 U357 ( .A(n112), .B(n109), .Y(n103) );
  OAI21X1 U358 ( .A0(n109), .A1(n113), .B0(n110), .Y(n104) );
  NAND2X1 U359 ( .A(n130), .B(n118), .Y(n116) );
  NOR2X1 U360 ( .A(n125), .B(n120), .Y(n118) );
  AOI21X1 U361 ( .A0(n172), .A1(n428), .B0(n169), .Y(n167) );
  NOR2X1 U362 ( .A(B[8]), .B(A[8]), .Y(n221) );
  NOR2X1 U363 ( .A(B[30]), .B(A[30]), .Y(n112) );
  NOR2X1 U364 ( .A(B[29]), .B(A[29]), .Y(n120) );
  INVX2 U365 ( .A(n115), .Y(n114) );
  AOI21X1 U366 ( .A0(n89), .A1(n104), .B0(n90), .Y(n84) );
  AOI21X2 U367 ( .A0(n115), .A1(n47), .B0(n48), .Y(n46) );
  OAI21X4 U368 ( .A0(n116), .A1(n144), .B0(n117), .Y(n115) );
  OAI21X2 U369 ( .A0(n173), .A1(n175), .B0(n174), .Y(n172) );
  AND2X4 U370 ( .A(n145), .B(n164), .Y(n426) );
  NOR2X4 U371 ( .A(n426), .B(n146), .Y(n144) );
  INVX1 U372 ( .A(n155), .Y(n153) );
  OR2XL U373 ( .A(B[24]), .B(A[24]), .Y(n429) );
  CLKINVXL U374 ( .A(n81), .Y(n79) );
  NAND2BX1 U375 ( .AN(n41), .B(n42), .Y(n1) );
  OAI21XL U376 ( .A0(n114), .A1(n65), .B0(n66), .Y(n64) );
  OAI21XL U377 ( .A0(n114), .A1(n101), .B0(n102), .Y(n100) );
  OAI21XL U378 ( .A0(n114), .A1(n56), .B0(n57), .Y(n55) );
  OAI21XL U379 ( .A0(n114), .A1(n76), .B0(n77), .Y(n75) );
  OAI21X1 U380 ( .A0(n73), .A1(n81), .B0(n74), .Y(n68) );
  NAND2BX1 U381 ( .AN(n120), .B(n121), .Y(n11) );
  OR2XL U382 ( .A(B[13]), .B(A[13]), .Y(n430) );
  OR2XL U383 ( .A(B[11]), .B(A[11]), .Y(n433) );
  NAND2X1 U384 ( .A(n89), .B(n103), .Y(n83) );
  CLKINVXL U385 ( .A(n84), .Y(n86) );
  AOI21XL U386 ( .A0(n86), .A1(n67), .B0(n68), .Y(n66) );
  CLKINVXL U387 ( .A(n104), .Y(n102) );
  CLKINVXL U388 ( .A(n130), .Y(n132) );
  CLKINVXL U389 ( .A(n184), .Y(n183) );
  CLKINVXL U390 ( .A(n99), .Y(n97) );
  CLKINVXL U391 ( .A(n98), .Y(n96) );
  NAND2XL U392 ( .A(n96), .B(n99), .Y(n8) );
  OAI21XL U393 ( .A0(n133), .A1(n125), .B0(n128), .Y(n124) );
  CLKINVX2 U394 ( .A(n158), .Y(n160) );
  CLKINVX2 U395 ( .A(n157), .Y(n273) );
  OAI21XL U396 ( .A0(n53), .A1(n63), .B0(n54), .Y(n52) );
  INVX1 U397 ( .A(n232), .Y(n231) );
  CLKINVXL U398 ( .A(n141), .Y(n270) );
  CLKINVXL U399 ( .A(n80), .Y(n78) );
  NAND2XL U400 ( .A(n428), .B(n171), .Y(n19) );
  NAND2BXL U401 ( .AN(n178), .B(n179), .Y(n21) );
  NAND2XL U402 ( .A(n273), .B(n158), .Y(n17) );
  NAND2BXL U403 ( .AN(n181), .B(n182), .Y(n22) );
  OAI21XL U404 ( .A0(n195), .A1(n193), .B0(n194), .Y(n192) );
  NAND2BXL U405 ( .AN(n193), .B(n194), .Y(n25) );
  NAND2XL U406 ( .A(n431), .B(n219), .Y(n31) );
  NAND2XL U407 ( .A(n432), .B(n227), .Y(n33) );
  NAND2XL U408 ( .A(n435), .B(n239), .Y(n36) );
  NAND2XL U409 ( .A(B[26]), .B(A[26]), .Y(n142) );
  NAND2XL U410 ( .A(B[30]), .B(A[30]), .Y(n113) );
  NAND2XL U411 ( .A(B[13]), .B(A[13]), .Y(n203) );
  NAND2XL U412 ( .A(B[21]), .B(A[21]), .Y(n171) );
  NAND2XL U413 ( .A(B[11]), .B(A[11]), .Y(n211) );
  NAND2XL U414 ( .A(B[8]), .B(A[8]), .Y(n222) );
  NAND2XL U415 ( .A(B[34]), .B(A[34]), .Y(n81) );
  NAND2XL U416 ( .A(B[24]), .B(A[24]), .Y(n155) );
  NAND2XL U417 ( .A(B[7]), .B(A[7]), .Y(n227) );
  NAND2XL U418 ( .A(B[22]), .B(A[22]), .Y(n166) );
  NAND2XL U419 ( .A(B[10]), .B(A[10]), .Y(n214) );
  NAND2XL U420 ( .A(B[36]), .B(A[36]), .Y(n63) );
  NAND2XL U421 ( .A(B[6]), .B(A[6]), .Y(n230) );
  NAND2XL U422 ( .A(B[9]), .B(A[9]), .Y(n219) );
  NAND2XL U423 ( .A(B[4]), .B(A[4]), .Y(n239) );
  NAND2XL U424 ( .A(n437), .B(A[38]), .Y(n45) );
  NAND2XL U425 ( .A(B[3]), .B(A[3]), .Y(n242) );
  INVX2 U426 ( .A(n438), .Y(n437) );
  INVX2 U427 ( .A(B[38]), .Y(n438) );
  INVX2 U428 ( .A(n83), .Y(n85) );
  OAI21XL U429 ( .A0(n114), .A1(n83), .B0(n84), .Y(n82) );
  INVX2 U430 ( .A(n164), .Y(n163) );
  OAI21X1 U431 ( .A0(n163), .A1(n150), .B0(n151), .Y(n149) );
  OAI21X1 U432 ( .A0(n46), .A1(n44), .B0(n45), .Y(n43) );
  NOR2X1 U433 ( .A(n60), .B(n53), .Y(n51) );
  NAND2XL U434 ( .A(n58), .B(n85), .Y(n56) );
  NOR2X1 U435 ( .A(n69), .B(n60), .Y(n58) );
  OAI21XL U436 ( .A0(n70), .A1(n60), .B0(n63), .Y(n59) );
  CLKINVXL U437 ( .A(n68), .Y(n70) );
  OAI21XL U438 ( .A0(n91), .A1(n99), .B0(n92), .Y(n90) );
  NOR2X1 U439 ( .A(n141), .B(n136), .Y(n130) );
  AOI21X1 U440 ( .A0(n131), .A1(n118), .B0(n119), .Y(n117) );
  OAI21X1 U441 ( .A0(n120), .A1(n128), .B0(n121), .Y(n119) );
  OAI21XL U442 ( .A0(n114), .A1(n94), .B0(n95), .Y(n93) );
  NAND2XL U443 ( .A(n103), .B(n96), .Y(n94) );
  OAI21XL U444 ( .A0(n114), .A1(n112), .B0(n113), .Y(n111) );
  NAND2XL U445 ( .A(n85), .B(n78), .Y(n76) );
  OAI21X1 U446 ( .A0(n142), .A1(n136), .B0(n137), .Y(n131) );
  INVX2 U447 ( .A(n171), .Y(n169) );
  NOR2X1 U448 ( .A(n150), .B(n147), .Y(n145) );
  AOI21X1 U449 ( .A0(n176), .A1(n184), .B0(n177), .Y(n175) );
  OAI21X1 U450 ( .A0(n178), .A1(n182), .B0(n179), .Y(n177) );
  NOR2X1 U451 ( .A(n181), .B(n178), .Y(n176) );
  AOI21XL U452 ( .A0(n123), .A1(n143), .B0(n124), .Y(n122) );
  NOR2X1 U453 ( .A(n132), .B(n125), .Y(n123) );
  CLKINVXL U454 ( .A(n131), .Y(n133) );
  AOI21XL U455 ( .A0(n143), .A1(n270), .B0(n140), .Y(n138) );
  INVX2 U456 ( .A(n142), .Y(n140) );
  OAI21X1 U457 ( .A0(n187), .A1(n185), .B0(n186), .Y(n184) );
  AOI21X1 U458 ( .A0(n188), .A1(n196), .B0(n189), .Y(n187) );
  OAI21X1 U459 ( .A0(n190), .A1(n194), .B0(n191), .Y(n189) );
  NOR2X1 U460 ( .A(n193), .B(n190), .Y(n188) );
  OAI21X1 U461 ( .A0(n199), .A1(n197), .B0(n198), .Y(n196) );
  INVX2 U462 ( .A(n203), .Y(n201) );
  INVX2 U463 ( .A(n211), .Y(n209) );
  OAI21X1 U464 ( .A0(n205), .A1(n207), .B0(n206), .Y(n204) );
  OAI21X1 U465 ( .A0(n213), .A1(n215), .B0(n214), .Y(n212) );
  AOI21X1 U466 ( .A0(n220), .A1(n431), .B0(n217), .Y(n215) );
  INVX2 U467 ( .A(n219), .Y(n217) );
  AOI21X1 U468 ( .A0(n228), .A1(n432), .B0(n225), .Y(n223) );
  INVX2 U469 ( .A(n227), .Y(n225) );
  OAI21X1 U470 ( .A0(n221), .A1(n223), .B0(n222), .Y(n220) );
  OAI21X1 U471 ( .A0(n241), .A1(n243), .B0(n242), .Y(n240) );
  INVX2 U472 ( .A(n247), .Y(n245) );
  OAI21X1 U473 ( .A0(n229), .A1(n231), .B0(n230), .Y(n228) );
  AOI21X1 U474 ( .A0(n435), .A1(n240), .B0(n237), .Y(n235) );
  INVX2 U475 ( .A(n239), .Y(n237) );
  OAI21X1 U476 ( .A0(n233), .A1(n235), .B0(n234), .Y(n232) );
  OAI2BB1X1 U477 ( .A0N(n436), .A1N(n254), .B0(n253), .Y(n427) );
  NAND2BX1 U478 ( .AN(n44), .B(n45), .Y(n2) );
  NAND2BX1 U479 ( .AN(n73), .B(n74), .Y(n5) );
  OAI21X1 U480 ( .A0(n163), .A1(n157), .B0(n158), .Y(n156) );
  NAND2BX1 U481 ( .AN(n53), .B(n54), .Y(n3) );
  NAND2X1 U482 ( .A(n273), .B(n429), .Y(n150) );
  NAND2BX1 U483 ( .AN(n60), .B(n63), .Y(n4) );
  NAND2XL U484 ( .A(n78), .B(n81), .Y(n6) );
  NAND2BX1 U485 ( .AN(n136), .B(n137), .Y(n13) );
  NAND2BX1 U486 ( .AN(n91), .B(n92), .Y(n7) );
  NAND2BX1 U487 ( .AN(n112), .B(n113), .Y(n10) );
  INVX2 U488 ( .A(n256), .Y(n254) );
  NAND2BX1 U489 ( .AN(n147), .B(n148), .Y(n15) );
  NAND2X1 U490 ( .A(n270), .B(n142), .Y(n14) );
  NAND2BX1 U491 ( .AN(n109), .B(n110), .Y(n9) );
  NAND2BX1 U492 ( .AN(n125), .B(n128), .Y(n12) );
  NAND2BX1 U493 ( .AN(n173), .B(n174), .Y(n20) );
  NAND2X1 U494 ( .A(n429), .B(n155), .Y(n16) );
  NAND2BX1 U495 ( .AN(n165), .B(n166), .Y(n18) );
  OAI21XL U496 ( .A0(n183), .A1(n181), .B0(n182), .Y(n180) );
  NAND2BX1 U497 ( .AN(n185), .B(n186), .Y(n23) );
  NAND2BX1 U498 ( .AN(n197), .B(n198), .Y(n26) );
  NAND2BX1 U499 ( .AN(n190), .B(n191), .Y(n24) );
  NAND2X1 U500 ( .A(n430), .B(n203), .Y(n27) );
  NAND2BX1 U501 ( .AN(n205), .B(n206), .Y(n28) );
  NAND2X1 U502 ( .A(n433), .B(n211), .Y(n29) );
  NAND2BX1 U503 ( .AN(n213), .B(n214), .Y(n30) );
  NAND2BX1 U504 ( .AN(n221), .B(n222), .Y(n32) );
  NAND2BX1 U505 ( .AN(n229), .B(n230), .Y(n34) );
  NAND2BX1 U506 ( .AN(n233), .B(n234), .Y(n35) );
  NAND2BX1 U507 ( .AN(n241), .B(n242), .Y(n37) );
  NAND2X1 U508 ( .A(n434), .B(n247), .Y(n38) );
  NAND2X1 U509 ( .A(n436), .B(n253), .Y(n39) );
  XNOR2X1 U510 ( .A(n43), .B(n1), .Y(SUM[39]) );
  NOR2X1 U511 ( .A(B[35]), .B(A[35]), .Y(n73) );
  XOR2X1 U512 ( .A(n46), .B(n2), .Y(SUM[38]) );
  XNOR2X1 U513 ( .A(n55), .B(n3), .Y(SUM[37]) );
  NAND2XL U514 ( .A(B[35]), .B(A[35]), .Y(n74) );
  NAND2XL U515 ( .A(B[37]), .B(A[37]), .Y(n54) );
  XNOR2X1 U516 ( .A(n64), .B(n4), .Y(SUM[36]) );
  XNOR2X1 U517 ( .A(n100), .B(n8), .Y(SUM[32]) );
  XNOR2X1 U518 ( .A(n111), .B(n9), .Y(SUM[31]) );
  XNOR2X1 U519 ( .A(n93), .B(n7), .Y(SUM[33]) );
  XNOR2X1 U520 ( .A(n82), .B(n6), .Y(SUM[34]) );
  XNOR2X1 U521 ( .A(n75), .B(n5), .Y(SUM[35]) );
  NOR2X1 U522 ( .A(B[20]), .B(A[20]), .Y(n173) );
  NOR2X1 U523 ( .A(B[32]), .B(A[32]), .Y(n98) );
  XOR2X1 U524 ( .A(n122), .B(n11), .Y(SUM[29]) );
  NOR2X1 U525 ( .A(B[26]), .B(A[26]), .Y(n141) );
  XOR2X1 U526 ( .A(n138), .B(n13), .Y(SUM[27]) );
  OR2X1 U527 ( .A(B[21]), .B(A[21]), .Y(n428) );
  NOR2X1 U528 ( .A(B[14]), .B(A[14]), .Y(n197) );
  NAND2X1 U529 ( .A(B[18]), .B(A[18]), .Y(n182) );
  NOR2X1 U530 ( .A(B[25]), .B(A[25]), .Y(n147) );
  NOR2X1 U531 ( .A(B[15]), .B(A[15]), .Y(n193) );
  XOR2X1 U532 ( .A(n114), .B(n10), .Y(SUM[30]) );
  NOR2X1 U533 ( .A(B[16]), .B(A[16]), .Y(n190) );
  NOR2X1 U534 ( .A(B[10]), .B(A[10]), .Y(n213) );
  OR2X1 U535 ( .A(B[9]), .B(A[9]), .Y(n431) );
  OR2X1 U536 ( .A(B[7]), .B(A[7]), .Y(n432) );
  NOR2X1 U537 ( .A(B[17]), .B(A[17]), .Y(n185) );
  NAND2XL U538 ( .A(B[20]), .B(A[20]), .Y(n174) );
  NAND2X1 U539 ( .A(B[23]), .B(A[23]), .Y(n158) );
  NOR2X1 U540 ( .A(B[28]), .B(A[28]), .Y(n125) );
  OR2XL U541 ( .A(B[2]), .B(A[2]), .Y(n434) );
  NOR2X1 U542 ( .A(B[12]), .B(A[12]), .Y(n205) );
  OR2X1 U543 ( .A(B[4]), .B(A[4]), .Y(n435) );
  NAND2XL U544 ( .A(B[19]), .B(A[19]), .Y(n179) );
  NAND2X1 U545 ( .A(B[32]), .B(A[32]), .Y(n99) );
  XNOR2X1 U546 ( .A(n143), .B(n14), .Y(SUM[26]) );
  NOR2X1 U547 ( .A(B[5]), .B(A[5]), .Y(n233) );
  NOR2X1 U548 ( .A(B[6]), .B(A[6]), .Y(n229) );
  NOR2X1 U549 ( .A(n437), .B(A[38]), .Y(n44) );
  NAND2X1 U550 ( .A(B[15]), .B(A[15]), .Y(n194) );
  OR2X1 U551 ( .A(B[1]), .B(A[1]), .Y(n436) );
  NAND2XL U552 ( .A(B[27]), .B(A[27]), .Y(n137) );
  NAND2XL U553 ( .A(B[14]), .B(A[14]), .Y(n198) );
  NAND2XL U554 ( .A(B[31]), .B(A[31]), .Y(n110) );
  NAND2XL U555 ( .A(B[28]), .B(A[28]), .Y(n128) );
  NAND2X1 U556 ( .A(n437), .B(A[39]), .Y(n42) );
  NOR2X1 U557 ( .A(n437), .B(A[39]), .Y(n41) );
  NAND2XL U558 ( .A(B[2]), .B(A[2]), .Y(n247) );
  NAND2XL U559 ( .A(B[33]), .B(A[33]), .Y(n92) );
  NAND2XL U560 ( .A(B[16]), .B(A[16]), .Y(n191) );
  XNOR2X1 U561 ( .A(n156), .B(n16), .Y(SUM[24]) );
  NOR2X1 U562 ( .A(B[3]), .B(A[3]), .Y(n241) );
  XNOR2X1 U563 ( .A(n149), .B(n15), .Y(SUM[25]) );
  NAND2XL U564 ( .A(B[17]), .B(A[17]), .Y(n186) );
  NAND2XL U565 ( .A(B[12]), .B(A[12]), .Y(n206) );
  NAND2XL U566 ( .A(B[29]), .B(A[29]), .Y(n121) );
  NAND2X1 U567 ( .A(B[1]), .B(A[1]), .Y(n253) );
  NOR2X1 U568 ( .A(B[23]), .B(A[23]), .Y(n157) );
  NAND2XL U569 ( .A(B[5]), .B(A[5]), .Y(n234) );
  NAND2XL U570 ( .A(B[25]), .B(A[25]), .Y(n148) );
  XOR2X1 U571 ( .A(n163), .B(n17), .Y(SUM[23]) );
  NOR2X1 U572 ( .A(B[22]), .B(A[22]), .Y(n165) );
  NAND2X1 U573 ( .A(B[0]), .B(A[0]), .Y(n256) );
  XNOR2X1 U574 ( .A(n172), .B(n19), .Y(SUM[21]) );
  XNOR2X1 U575 ( .A(n192), .B(n24), .Y(SUM[16]) );
  XNOR2X1 U576 ( .A(n180), .B(n21), .Y(SUM[19]) );
  XOR2X1 U577 ( .A(n25), .B(n195), .Y(SUM[15]) );
  XOR2X1 U578 ( .A(n183), .B(n22), .Y(SUM[18]) );
  XNOR2XL U579 ( .A(n27), .B(n204), .Y(SUM[13]) );
  XNOR2XL U580 ( .A(n29), .B(n212), .Y(SUM[11]) );
  XOR2XL U581 ( .A(n30), .B(n215), .Y(SUM[10]) );
  XNOR2XL U582 ( .A(n31), .B(n220), .Y(SUM[9]) );
  XOR2XL U583 ( .A(n32), .B(n223), .Y(SUM[8]) );
  XNOR2XL U584 ( .A(n33), .B(n228), .Y(SUM[7]) );
  XOR2XL U585 ( .A(n34), .B(n231), .Y(SUM[6]) );
  XNOR2XL U586 ( .A(n36), .B(n240), .Y(SUM[4]) );
  XNOR2X1 U587 ( .A(n38), .B(n427), .Y(SUM[2]) );
  XNOR2X1 U588 ( .A(n39), .B(n254), .Y(SUM[1]) );
  NAND2BX1 U589 ( .AN(n255), .B(n256), .Y(n40) );
  NOR2X1 U590 ( .A(B[0]), .B(A[0]), .Y(n255) );
  INVX2 U591 ( .A(n40), .Y(SUM[0]) );
  CLKINVXL U592 ( .A(n196), .Y(n195) );
  XOR2X1 U593 ( .A(n28), .B(n207), .Y(SUM[12]) );
  NAND2XL U594 ( .A(n85), .B(n67), .Y(n65) );
  NAND2X1 U595 ( .A(n67), .B(n51), .Y(n49) );
  INVX2 U596 ( .A(n103), .Y(n101) );
  XOR2X1 U597 ( .A(n187), .B(n23), .Y(SUM[17]) );
  NOR2X1 U598 ( .A(n49), .B(n83), .Y(n47) );
  XOR2X1 U599 ( .A(n129), .B(n12), .Y(SUM[28]) );
  INVX1 U600 ( .A(n144), .Y(n143) );
  XOR2XL U601 ( .A(n18), .B(n167), .Y(SUM[22]) );
  XOR2XL U602 ( .A(n35), .B(n235), .Y(SUM[5]) );
  XOR2XL U603 ( .A(n37), .B(n243), .Y(SUM[3]) );
  XOR2XL U604 ( .A(n20), .B(n175), .Y(SUM[20]) );
  XOR2XL U605 ( .A(n26), .B(n199), .Y(SUM[14]) );
endmodule


module MMSA_DW01_add_40 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n63, n64, n65, n66, n67, n68, n69, n70, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n128, n129, n130, n131, n132, n133,
         n136, n137, n138, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n153, n155, n156, n157, n158, n160, n163,
         n164, n165, n166, n167, n169, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n201, n203, n204, n205, n206, n207, n209, n211, n212, n213,
         n214, n215, n217, n219, n220, n221, n222, n223, n225, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n237, n239, n240, n241,
         n242, n243, n245, n247, n253, n254, n255, n256, n270, n273, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435;

  AOI21X1 U13 ( .A0(n115), .A1(n47), .B0(n48), .Y(n46) );
  AOI21X1 U17 ( .A0(n51), .A1(n68), .B0(n52), .Y(n50) );
  AOI21X1 U27 ( .A0(n58), .A1(n86), .B0(n59), .Y(n57) );
  AOI21X1 U53 ( .A0(n86), .A1(n78), .B0(n79), .Y(n77) );
  AOI21X1 U77 ( .A0(n104), .A1(n96), .B0(n97), .Y(n95) );
  AOI21X1 U108 ( .A0(n131), .A1(n118), .B0(n119), .Y(n117) );
  AOI21X1 U116 ( .A0(n123), .A1(n143), .B0(n124), .Y(n122) );
  AOI21X1 U138 ( .A0(n143), .A1(n270), .B0(n140), .Y(n138) );
  AOI21X1 U157 ( .A0(n426), .A1(n160), .B0(n153), .Y(n151) );
  AOI21X1 U266 ( .A0(n220), .A1(n431), .B0(n217), .Y(n215) );
  AOI21X1 U315 ( .A0(n432), .A1(n424), .B0(n245), .Y(n243) );
  NOR2X2 U340 ( .A(B[31]), .B(A[31]), .Y(n109) );
  OAI21X2 U341 ( .A0(n109), .A1(n113), .B0(n110), .Y(n104) );
  NOR2X1 U342 ( .A(B[34]), .B(A[34]), .Y(n80) );
  NOR2X2 U343 ( .A(B[33]), .B(A[33]), .Y(n91) );
  NAND2X1 U344 ( .A(n89), .B(n103), .Y(n83) );
  NOR2X2 U345 ( .A(n91), .B(n98), .Y(n89) );
  OAI21X2 U346 ( .A0(n73), .A1(n81), .B0(n74), .Y(n68) );
  NOR2X2 U347 ( .A(B[35]), .B(A[35]), .Y(n73) );
  OAI21X2 U348 ( .A0(n187), .A1(n185), .B0(n186), .Y(n184) );
  AOI21X2 U349 ( .A0(n188), .A1(n196), .B0(n189), .Y(n187) );
  NOR2X2 U350 ( .A(n80), .B(n73), .Y(n67) );
  NOR2X1 U351 ( .A(B[18]), .B(A[18]), .Y(n181) );
  OAI21X1 U352 ( .A0(n199), .A1(n197), .B0(n198), .Y(n196) );
  NOR2X1 U353 ( .A(n112), .B(n109), .Y(n103) );
  NOR2X1 U354 ( .A(n125), .B(n120), .Y(n118) );
  NOR2X1 U355 ( .A(B[25]), .B(A[25]), .Y(n147) );
  OAI21X1 U356 ( .A0(n173), .A1(n175), .B0(n174), .Y(n172) );
  NOR2X1 U357 ( .A(B[28]), .B(A[28]), .Y(n125) );
  NOR2X1 U358 ( .A(B[30]), .B(A[30]), .Y(n112) );
  NOR2X1 U359 ( .A(B[27]), .B(A[27]), .Y(n136) );
  OAI21X1 U360 ( .A0(n151), .A1(n147), .B0(n148), .Y(n146) );
  OAI21X2 U361 ( .A0(n165), .A1(n167), .B0(n166), .Y(n164) );
  OAI21X2 U362 ( .A0(n116), .A1(n144), .B0(n117), .Y(n115) );
  AOI21X2 U363 ( .A0(n145), .A1(n164), .B0(n146), .Y(n144) );
  AOI21XL U364 ( .A0(n89), .A1(n104), .B0(n90), .Y(n423) );
  AOI21XL U365 ( .A0(n89), .A1(n104), .B0(n90), .Y(n84) );
  AOI21XL U366 ( .A0(n86), .A1(n67), .B0(n68), .Y(n66) );
  OAI21XL U367 ( .A0(n114), .A1(n65), .B0(n66), .Y(n64) );
  OAI21XL U368 ( .A0(n114), .A1(n56), .B0(n57), .Y(n55) );
  OAI21X1 U369 ( .A0(n91), .A1(n99), .B0(n92), .Y(n90) );
  NAND2XL U370 ( .A(n58), .B(n85), .Y(n56) );
  CLKINVXL U371 ( .A(n81), .Y(n79) );
  OAI21XL U372 ( .A0(n53), .A1(n63), .B0(n54), .Y(n52) );
  NAND2BX1 U373 ( .AN(n41), .B(n42), .Y(n1) );
  OAI21XL U374 ( .A0(n114), .A1(n76), .B0(n77), .Y(n75) );
  NOR2X1 U375 ( .A(B[36]), .B(A[36]), .Y(n60) );
  XNOR2XL U376 ( .A(n36), .B(n240), .Y(SUM[4]) );
  XNOR2XL U377 ( .A(n38), .B(n424), .Y(SUM[2]) );
  CLKINVXL U378 ( .A(n104), .Y(n102) );
  OAI21XL U379 ( .A0(n163), .A1(n150), .B0(n151), .Y(n149) );
  CLKINVXL U380 ( .A(n130), .Y(n132) );
  CLKINVXL U381 ( .A(n184), .Y(n183) );
  OAI21X1 U382 ( .A0(n46), .A1(n44), .B0(n45), .Y(n43) );
  CLKINVXL U383 ( .A(n99), .Y(n97) );
  CLKINVXL U384 ( .A(n98), .Y(n96) );
  CLKINVX1 U385 ( .A(n219), .Y(n217) );
  NAND2XL U386 ( .A(n96), .B(n99), .Y(n8) );
  CLKINVX2 U387 ( .A(n157), .Y(n273) );
  OAI21XL U388 ( .A0(n163), .A1(n157), .B0(n158), .Y(n156) );
  CLKINVX1 U389 ( .A(n227), .Y(n225) );
  INVX1 U390 ( .A(n232), .Y(n231) );
  CLKINVXL U391 ( .A(n141), .Y(n270) );
  CLKINVXL U392 ( .A(n80), .Y(n78) );
  NAND2BXL U393 ( .AN(n125), .B(n128), .Y(n12) );
  OAI21XL U394 ( .A0(n195), .A1(n193), .B0(n194), .Y(n192) );
  NAND2XL U395 ( .A(n429), .B(n211), .Y(n29) );
  NAND2XL U396 ( .A(n431), .B(n219), .Y(n31) );
  NAND2XL U397 ( .A(n430), .B(n227), .Y(n33) );
  OR2XL U398 ( .A(B[24]), .B(A[24]), .Y(n426) );
  NAND2XL U399 ( .A(B[24]), .B(A[24]), .Y(n155) );
  NAND2XL U400 ( .A(B[27]), .B(A[27]), .Y(n137) );
  NAND2XL U401 ( .A(B[30]), .B(A[30]), .Y(n113) );
  NAND2XL U402 ( .A(B[26]), .B(A[26]), .Y(n142) );
  NAND2XL U403 ( .A(B[18]), .B(A[18]), .Y(n182) );
  NAND2XL U404 ( .A(B[15]), .B(A[15]), .Y(n194) );
  NAND2XL U405 ( .A(B[8]), .B(A[8]), .Y(n222) );
  OR2XL U406 ( .A(B[13]), .B(A[13]), .Y(n427) );
  NAND2XL U407 ( .A(B[13]), .B(A[13]), .Y(n203) );
  NAND2XL U408 ( .A(B[23]), .B(A[23]), .Y(n158) );
  OR2XL U409 ( .A(B[21]), .B(A[21]), .Y(n425) );
  NAND2XL U410 ( .A(B[21]), .B(A[21]), .Y(n171) );
  OR2XL U411 ( .A(B[7]), .B(A[7]), .Y(n430) );
  NAND2XL U412 ( .A(B[14]), .B(A[14]), .Y(n198) );
  NAND2XL U413 ( .A(B[34]), .B(A[34]), .Y(n81) );
  NAND2XL U414 ( .A(B[36]), .B(A[36]), .Y(n63) );
  NAND2XL U415 ( .A(B[22]), .B(A[22]), .Y(n166) );
  NAND2XL U416 ( .A(n434), .B(A[38]), .Y(n45) );
  INVX2 U417 ( .A(n435), .Y(n434) );
  INVX2 U418 ( .A(B[38]), .Y(n435) );
  INVX2 U419 ( .A(n83), .Y(n85) );
  NOR2X1 U420 ( .A(n49), .B(n83), .Y(n47) );
  OAI21X1 U421 ( .A0(n84), .A1(n49), .B0(n50), .Y(n48) );
  NAND2X1 U422 ( .A(n67), .B(n51), .Y(n49) );
  INVX2 U423 ( .A(n67), .Y(n69) );
  INVX2 U424 ( .A(n115), .Y(n114) );
  INVX2 U425 ( .A(n144), .Y(n143) );
  OAI21XL U426 ( .A0(n114), .A1(n101), .B0(n102), .Y(n100) );
  CLKINVXL U427 ( .A(n103), .Y(n101) );
  INVX2 U428 ( .A(n164), .Y(n163) );
  INVX2 U429 ( .A(n196), .Y(n195) );
  NOR2X1 U430 ( .A(n60), .B(n53), .Y(n51) );
  OAI21X1 U431 ( .A0(n70), .A1(n60), .B0(n63), .Y(n59) );
  CLKINVXL U432 ( .A(n68), .Y(n70) );
  NAND2XL U433 ( .A(n85), .B(n78), .Y(n76) );
  OAI21X1 U434 ( .A0(n142), .A1(n136), .B0(n137), .Y(n131) );
  NAND2X1 U435 ( .A(n130), .B(n118), .Y(n116) );
  OAI21X1 U436 ( .A0(n190), .A1(n194), .B0(n191), .Y(n189) );
  NOR2X1 U437 ( .A(n193), .B(n190), .Y(n188) );
  NOR2X1 U438 ( .A(n150), .B(n147), .Y(n145) );
  AOI21X1 U439 ( .A0(n176), .A1(n184), .B0(n177), .Y(n175) );
  OAI21X1 U440 ( .A0(n178), .A1(n182), .B0(n179), .Y(n177) );
  NOR2X1 U441 ( .A(n181), .B(n178), .Y(n176) );
  AOI21X1 U442 ( .A0(n172), .A1(n425), .B0(n169), .Y(n167) );
  INVX2 U443 ( .A(n171), .Y(n169) );
  AOI21X1 U444 ( .A0(n204), .A1(n427), .B0(n201), .Y(n199) );
  INVX2 U445 ( .A(n203), .Y(n201) );
  AOI21X1 U446 ( .A0(n228), .A1(n430), .B0(n225), .Y(n223) );
  OAI21X1 U447 ( .A0(n205), .A1(n207), .B0(n206), .Y(n204) );
  OAI21X1 U448 ( .A0(n213), .A1(n215), .B0(n214), .Y(n212) );
  OAI21X1 U449 ( .A0(n229), .A1(n231), .B0(n230), .Y(n228) );
  AOI21X1 U450 ( .A0(n428), .A1(n240), .B0(n237), .Y(n235) );
  INVX2 U451 ( .A(n239), .Y(n237) );
  OAI21X1 U452 ( .A0(n221), .A1(n223), .B0(n222), .Y(n220) );
  AOI21X1 U453 ( .A0(n429), .A1(n212), .B0(n209), .Y(n207) );
  INVX2 U454 ( .A(n211), .Y(n209) );
  OAI21X1 U455 ( .A0(n233), .A1(n235), .B0(n234), .Y(n232) );
  NOR2X1 U456 ( .A(n141), .B(n136), .Y(n130) );
  INVX2 U457 ( .A(n155), .Y(n153) );
  INVX2 U458 ( .A(n158), .Y(n160) );
  OAI21XL U459 ( .A0(n114), .A1(n112), .B0(n113), .Y(n111) );
  OAI21XL U460 ( .A0(n114), .A1(n94), .B0(n95), .Y(n93) );
  NAND2XL U461 ( .A(n103), .B(n96), .Y(n94) );
  OAI21XL U462 ( .A0(n133), .A1(n125), .B0(n128), .Y(n124) );
  NOR2X1 U463 ( .A(n132), .B(n125), .Y(n123) );
  CLKINVXL U464 ( .A(n131), .Y(n133) );
  NAND2X1 U465 ( .A(n273), .B(n426), .Y(n150) );
  INVX2 U466 ( .A(n142), .Y(n140) );
  NAND2BX1 U467 ( .AN(n44), .B(n45), .Y(n2) );
  NAND2BX1 U468 ( .AN(n73), .B(n74), .Y(n5) );
  INVX2 U469 ( .A(n247), .Y(n245) );
  OAI21X1 U470 ( .A0(n241), .A1(n243), .B0(n242), .Y(n240) );
  NAND2XL U471 ( .A(n78), .B(n81), .Y(n6) );
  NAND2BX1 U472 ( .AN(n53), .B(n54), .Y(n3) );
  NAND2BX1 U473 ( .AN(n60), .B(n63), .Y(n4) );
  OAI2BB1X1 U474 ( .A0N(n433), .A1N(n254), .B0(n253), .Y(n424) );
  NAND2BX1 U475 ( .AN(n136), .B(n137), .Y(n13) );
  NAND2BX1 U476 ( .AN(n120), .B(n121), .Y(n11) );
  NAND2BX1 U477 ( .AN(n91), .B(n92), .Y(n7) );
  NAND2BX1 U478 ( .AN(n112), .B(n113), .Y(n10) );
  NAND2BX1 U479 ( .AN(n147), .B(n148), .Y(n15) );
  NAND2BX1 U480 ( .AN(n109), .B(n110), .Y(n9) );
  NAND2X1 U481 ( .A(n270), .B(n142), .Y(n14) );
  INVX2 U482 ( .A(n256), .Y(n254) );
  NAND2XL U483 ( .A(n273), .B(n158), .Y(n17) );
  NAND2BX1 U484 ( .AN(n173), .B(n174), .Y(n20) );
  NAND2X1 U485 ( .A(n425), .B(n171), .Y(n19) );
  OAI21XL U486 ( .A0(n183), .A1(n181), .B0(n182), .Y(n180) );
  NAND2BX1 U487 ( .AN(n165), .B(n166), .Y(n18) );
  NAND2X1 U488 ( .A(n426), .B(n155), .Y(n16) );
  NAND2BX1 U489 ( .AN(n178), .B(n179), .Y(n21) );
  NAND2BX1 U490 ( .AN(n181), .B(n182), .Y(n22) );
  NAND2BX1 U491 ( .AN(n185), .B(n186), .Y(n23) );
  NAND2BX1 U492 ( .AN(n197), .B(n198), .Y(n26) );
  NAND2BX1 U493 ( .AN(n190), .B(n191), .Y(n24) );
  NAND2BX1 U494 ( .AN(n193), .B(n194), .Y(n25) );
  NAND2X1 U495 ( .A(n427), .B(n203), .Y(n27) );
  NAND2BX1 U496 ( .AN(n205), .B(n206), .Y(n28) );
  NAND2BX1 U497 ( .AN(n213), .B(n214), .Y(n30) );
  NAND2BX1 U498 ( .AN(n221), .B(n222), .Y(n32) );
  NAND2BX1 U499 ( .AN(n229), .B(n230), .Y(n34) );
  NAND2BX1 U500 ( .AN(n233), .B(n234), .Y(n35) );
  NAND2XL U501 ( .A(n428), .B(n239), .Y(n36) );
  NAND2BX1 U502 ( .AN(n241), .B(n242), .Y(n37) );
  NAND2X1 U503 ( .A(n432), .B(n247), .Y(n38) );
  NAND2X1 U504 ( .A(n433), .B(n253), .Y(n39) );
  XNOR2X1 U505 ( .A(n43), .B(n1), .Y(SUM[39]) );
  NOR2X1 U506 ( .A(B[37]), .B(A[37]), .Y(n53) );
  XNOR2X1 U507 ( .A(n55), .B(n3), .Y(SUM[37]) );
  NAND2XL U508 ( .A(B[35]), .B(A[35]), .Y(n74) );
  NAND2XL U509 ( .A(B[37]), .B(A[37]), .Y(n54) );
  XNOR2X1 U510 ( .A(n64), .B(n4), .Y(SUM[36]) );
  XNOR2X1 U511 ( .A(n75), .B(n5), .Y(SUM[35]) );
  NOR2X1 U512 ( .A(B[16]), .B(A[16]), .Y(n190) );
  NOR2X1 U513 ( .A(B[20]), .B(A[20]), .Y(n173) );
  NOR2X1 U514 ( .A(B[14]), .B(A[14]), .Y(n197) );
  NOR2X1 U515 ( .A(B[29]), .B(A[29]), .Y(n120) );
  NOR2X1 U516 ( .A(B[19]), .B(A[19]), .Y(n178) );
  NOR2X1 U517 ( .A(B[12]), .B(A[12]), .Y(n205) );
  NAND2XL U518 ( .A(B[28]), .B(A[28]), .Y(n128) );
  NOR2X1 U519 ( .A(B[26]), .B(A[26]), .Y(n141) );
  NOR2X1 U520 ( .A(B[15]), .B(A[15]), .Y(n193) );
  NOR2X1 U521 ( .A(B[32]), .B(A[32]), .Y(n98) );
  XOR2X1 U522 ( .A(n129), .B(n12), .Y(SUM[28]) );
  NOR2X1 U523 ( .A(B[17]), .B(A[17]), .Y(n185) );
  OR2XL U524 ( .A(B[4]), .B(A[4]), .Y(n428) );
  XNOR2X1 U525 ( .A(n111), .B(n9), .Y(SUM[31]) );
  NAND2XL U526 ( .A(B[20]), .B(A[20]), .Y(n174) );
  XNOR2X1 U527 ( .A(n100), .B(n8), .Y(SUM[32]) );
  XNOR2X1 U528 ( .A(n93), .B(n7), .Y(SUM[33]) );
  NAND2XL U529 ( .A(B[29]), .B(A[29]), .Y(n121) );
  XOR2X1 U530 ( .A(n122), .B(n11), .Y(SUM[29]) );
  NOR2X1 U531 ( .A(B[5]), .B(A[5]), .Y(n233) );
  NAND2XL U532 ( .A(B[19]), .B(A[19]), .Y(n179) );
  NOR2X1 U533 ( .A(B[23]), .B(A[23]), .Y(n157) );
  XOR2X1 U534 ( .A(n138), .B(n13), .Y(SUM[27]) );
  NAND2XL U535 ( .A(B[16]), .B(A[16]), .Y(n191) );
  NOR2X1 U536 ( .A(n434), .B(A[38]), .Y(n44) );
  NAND2XL U537 ( .A(B[12]), .B(A[12]), .Y(n206) );
  NAND2X1 U538 ( .A(B[32]), .B(A[32]), .Y(n99) );
  OR2XL U539 ( .A(B[11]), .B(A[11]), .Y(n429) );
  XOR2X1 U540 ( .A(n114), .B(n10), .Y(SUM[30]) );
  NOR2X1 U541 ( .A(B[10]), .B(A[10]), .Y(n213) );
  NOR2X1 U542 ( .A(B[6]), .B(A[6]), .Y(n229) );
  NAND2XL U543 ( .A(B[31]), .B(A[31]), .Y(n110) );
  NAND2XL U544 ( .A(B[25]), .B(A[25]), .Y(n148) );
  OR2XL U545 ( .A(B[9]), .B(A[9]), .Y(n431) );
  NAND2XL U546 ( .A(B[33]), .B(A[33]), .Y(n92) );
  NAND2XL U547 ( .A(B[11]), .B(A[11]), .Y(n211) );
  NAND2XL U548 ( .A(n434), .B(A[39]), .Y(n42) );
  NOR2X1 U549 ( .A(n434), .B(A[39]), .Y(n41) );
  NAND2XL U550 ( .A(B[17]), .B(A[17]), .Y(n186) );
  NAND2XL U551 ( .A(B[5]), .B(A[5]), .Y(n234) );
  OR2XL U552 ( .A(B[2]), .B(A[2]), .Y(n432) );
  NAND2XL U553 ( .A(B[7]), .B(A[7]), .Y(n227) );
  NAND2XL U554 ( .A(B[9]), .B(A[9]), .Y(n219) );
  NAND2XL U555 ( .A(B[10]), .B(A[10]), .Y(n214) );
  NOR2X1 U556 ( .A(B[8]), .B(A[8]), .Y(n221) );
  NOR2X1 U557 ( .A(B[3]), .B(A[3]), .Y(n241) );
  NAND2XL U558 ( .A(B[6]), .B(A[6]), .Y(n230) );
  NAND2XL U559 ( .A(B[2]), .B(A[2]), .Y(n247) );
  OR2XL U560 ( .A(B[1]), .B(A[1]), .Y(n433) );
  NOR2X1 U561 ( .A(B[22]), .B(A[22]), .Y(n165) );
  NAND2XL U562 ( .A(B[1]), .B(A[1]), .Y(n253) );
  NAND2XL U563 ( .A(B[3]), .B(A[3]), .Y(n242) );
  XNOR2X1 U564 ( .A(n143), .B(n14), .Y(SUM[26]) );
  XNOR2X1 U565 ( .A(n156), .B(n16), .Y(SUM[24]) );
  XNOR2X1 U566 ( .A(n149), .B(n15), .Y(SUM[25]) );
  XOR2X1 U567 ( .A(n163), .B(n17), .Y(SUM[23]) );
  NAND2X1 U568 ( .A(B[0]), .B(A[0]), .Y(n256) );
  XNOR2X1 U569 ( .A(n172), .B(n19), .Y(SUM[21]) );
  XNOR2X1 U570 ( .A(n180), .B(n21), .Y(SUM[19]) );
  XOR2X1 U571 ( .A(n183), .B(n22), .Y(SUM[18]) );
  XNOR2X1 U572 ( .A(n192), .B(n24), .Y(SUM[16]) );
  XOR2XL U573 ( .A(n26), .B(n199), .Y(SUM[14]) );
  XOR2X1 U574 ( .A(n25), .B(n195), .Y(SUM[15]) );
  XNOR2XL U575 ( .A(n27), .B(n204), .Y(SUM[13]) );
  XNOR2XL U576 ( .A(n31), .B(n220), .Y(SUM[9]) );
  XOR2XL U577 ( .A(n32), .B(n223), .Y(SUM[8]) );
  XNOR2XL U578 ( .A(n33), .B(n228), .Y(SUM[7]) );
  XOR2XL U579 ( .A(n34), .B(n231), .Y(SUM[6]) );
  XNOR2X1 U580 ( .A(n39), .B(n254), .Y(SUM[1]) );
  NAND2BX1 U581 ( .AN(n255), .B(n256), .Y(n40) );
  NOR2X1 U582 ( .A(B[0]), .B(A[0]), .Y(n255) );
  INVX2 U583 ( .A(n40), .Y(SUM[0]) );
  NAND2XL U584 ( .A(B[4]), .B(A[4]), .Y(n239) );
  AOI21XL U585 ( .A0(n143), .A1(n130), .B0(n131), .Y(n129) );
  XNOR2XL U586 ( .A(n29), .B(n212), .Y(SUM[11]) );
  XOR2XL U587 ( .A(n35), .B(n235), .Y(SUM[5]) );
  XOR2X1 U588 ( .A(n187), .B(n23), .Y(SUM[17]) );
  XOR2XL U589 ( .A(n37), .B(n243), .Y(SUM[3]) );
  NAND2XL U590 ( .A(n85), .B(n67), .Y(n65) );
  INVX2 U591 ( .A(n423), .Y(n86) );
  NOR2X1 U592 ( .A(n69), .B(n60), .Y(n58) );
  XNOR2X1 U593 ( .A(n82), .B(n6), .Y(SUM[34]) );
  OAI21XL U594 ( .A0(n120), .A1(n128), .B0(n121), .Y(n119) );
  XOR2XL U595 ( .A(n18), .B(n167), .Y(SUM[22]) );
  XOR2XL U596 ( .A(n20), .B(n175), .Y(SUM[20]) );
  XOR2XL U597 ( .A(n28), .B(n207), .Y(SUM[12]) );
  XOR2XL U598 ( .A(n30), .B(n215), .Y(SUM[10]) );
  XOR2X1 U599 ( .A(n46), .B(n2), .Y(SUM[38]) );
  OAI21XL U600 ( .A0(n114), .A1(n83), .B0(n423), .Y(n82) );
endmodule


module MMSA_DW01_add_39 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n63, n64, n65, n66, n67, n68, n69, n70, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n128, n129, n130, n131, n133, n136,
         n137, n138, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n153, n155, n156, n157, n158, n160, n163, n164,
         n165, n166, n167, n169, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n201, n203, n204, n205, n206, n207, n209, n211, n212, n213, n214,
         n215, n217, n219, n220, n221, n222, n223, n225, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n237, n239, n240, n241, n242,
         n243, n245, n247, n253, n254, n255, n256, n270, n273, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439;

  AOI21X1 U17 ( .A0(n51), .A1(n68), .B0(n52), .Y(n50) );
  AOI21X1 U27 ( .A0(n58), .A1(n86), .B0(n59), .Y(n57) );
  NOR2X2 U34 ( .A(B[36]), .B(A[36]), .Y(n60) );
  AOI21X1 U39 ( .A0(n86), .A1(n67), .B0(n68), .Y(n66) );
  NOR2X2 U44 ( .A(n80), .B(n73), .Y(n67) );
  NOR2X2 U48 ( .A(B[35]), .B(A[35]), .Y(n73) );
  AOI21X1 U53 ( .A0(n86), .A1(n78), .B0(n79), .Y(n77) );
  AOI21X1 U77 ( .A0(n104), .A1(n96), .B0(n97), .Y(n95) );
  AOI21X1 U126 ( .A0(n143), .A1(n130), .B0(n131), .Y(n129) );
  AOI21X1 U138 ( .A0(n143), .A1(n270), .B0(n140), .Y(n138) );
  AOI21X1 U157 ( .A0(n431), .A1(n160), .B0(n153), .Y(n151) );
  AOI21X1 U280 ( .A0(n228), .A1(n432), .B0(n225), .Y(n223) );
  NOR2X2 U340 ( .A(B[29]), .B(A[29]), .Y(n120) );
  NAND2X4 U341 ( .A(n425), .B(n117), .Y(n115) );
  OAI21X2 U342 ( .A0(n84), .A1(n49), .B0(n50), .Y(n48) );
  NOR2X1 U343 ( .A(B[34]), .B(A[34]), .Y(n80) );
  AOI21X2 U344 ( .A0(n115), .A1(n47), .B0(n48), .Y(n46) );
  NAND2X1 U345 ( .A(B[23]), .B(A[23]), .Y(n158) );
  NAND2X2 U346 ( .A(n423), .B(n424), .Y(n425) );
  INVX4 U347 ( .A(n116), .Y(n423) );
  INVX2 U348 ( .A(n427), .Y(n424) );
  AOI21X2 U349 ( .A0(n131), .A1(n118), .B0(n119), .Y(n117) );
  INVX1 U350 ( .A(n115), .Y(n114) );
  NOR2X1 U351 ( .A(n91), .B(n98), .Y(n89) );
  NOR2X1 U352 ( .A(n60), .B(n53), .Y(n51) );
  OAI21X1 U353 ( .A0(n91), .A1(n99), .B0(n92), .Y(n90) );
  NOR2X1 U354 ( .A(B[33]), .B(A[33]), .Y(n91) );
  NAND2X1 U355 ( .A(n67), .B(n51), .Y(n49) );
  OAI21X2 U356 ( .A0(n73), .A1(n81), .B0(n74), .Y(n68) );
  AOI21X1 U357 ( .A0(n89), .A1(n104), .B0(n90), .Y(n84) );
  NAND2X1 U358 ( .A(B[34]), .B(A[34]), .Y(n81) );
  NAND2XL U359 ( .A(B[26]), .B(A[26]), .Y(n142) );
  OAI21X1 U360 ( .A0(n165), .A1(n167), .B0(n166), .Y(n164) );
  BUFX1 U361 ( .A(n164), .Y(n426) );
  AOI21X1 U362 ( .A0(n145), .A1(n164), .B0(n146), .Y(n427) );
  CLKINVXL U363 ( .A(n155), .Y(n153) );
  AOI21XL U364 ( .A0(n145), .A1(n426), .B0(n146), .Y(n144) );
  CLKINVX2 U365 ( .A(n158), .Y(n160) );
  NAND2XL U366 ( .A(B[18]), .B(A[18]), .Y(n182) );
  NAND2XL U367 ( .A(B[15]), .B(A[15]), .Y(n194) );
  OR2XL U368 ( .A(B[24]), .B(A[24]), .Y(n431) );
  NAND2BX1 U369 ( .AN(n41), .B(n42), .Y(n1) );
  OR2XL U370 ( .A(B[4]), .B(A[4]), .Y(n433) );
  CLKINVXL U371 ( .A(n104), .Y(n102) );
  NAND2BX1 U372 ( .AN(n125), .B(n128), .Y(n12) );
  XNOR2XL U373 ( .A(n31), .B(n220), .Y(SUM[9]) );
  XOR2XL U374 ( .A(n35), .B(n235), .Y(SUM[5]) );
  XNOR2XL U375 ( .A(n36), .B(n240), .Y(SUM[4]) );
  XOR2XL U376 ( .A(n37), .B(n243), .Y(SUM[3]) );
  XNOR2XL U377 ( .A(n38), .B(n428), .Y(SUM[2]) );
  CLKINVXL U378 ( .A(n83), .Y(n85) );
  CLKINVXL U379 ( .A(n84), .Y(n86) );
  CLKINVXL U380 ( .A(n103), .Y(n101) );
  INVX1 U381 ( .A(n131), .Y(n133) );
  CLKINVXL U382 ( .A(n184), .Y(n183) );
  CLKINVXL U383 ( .A(n196), .Y(n195) );
  OAI21X1 U384 ( .A0(n120), .A1(n128), .B0(n121), .Y(n119) );
  OAI21X1 U385 ( .A0(n114), .A1(n56), .B0(n57), .Y(n55) );
  CLKINVXL U386 ( .A(n99), .Y(n97) );
  NOR2BXL U387 ( .AN(n130), .B(n125), .Y(n123) );
  OAI21X2 U388 ( .A0(n109), .A1(n113), .B0(n110), .Y(n104) );
  CLKINVXL U389 ( .A(n98), .Y(n96) );
  NAND2XL U390 ( .A(n96), .B(n99), .Y(n8) );
  CLKINVX2 U391 ( .A(n157), .Y(n273) );
  OAI21XL U392 ( .A0(n163), .A1(n157), .B0(n158), .Y(n156) );
  OAI21XL U393 ( .A0(n53), .A1(n63), .B0(n54), .Y(n52) );
  NAND2XL U394 ( .A(n431), .B(n155), .Y(n16) );
  INVX1 U395 ( .A(n232), .Y(n231) );
  CLKINVX1 U396 ( .A(n239), .Y(n237) );
  CLKINVXL U397 ( .A(n141), .Y(n270) );
  NAND2XL U398 ( .A(n273), .B(n158), .Y(n17) );
  NAND2XL U399 ( .A(n429), .B(n171), .Y(n19) );
  OAI21XL U400 ( .A0(n183), .A1(n181), .B0(n182), .Y(n180) );
  OAI21XL U401 ( .A0(n195), .A1(n193), .B0(n194), .Y(n192) );
  NAND2XL U402 ( .A(n430), .B(n203), .Y(n27) );
  NAND2XL U403 ( .A(n434), .B(n211), .Y(n29) );
  NAND2XL U404 ( .A(n436), .B(n219), .Y(n31) );
  NAND2XL U405 ( .A(n432), .B(n227), .Y(n33) );
  NAND2XL U406 ( .A(n433), .B(n239), .Y(n36) );
  NAND2XL U407 ( .A(B[30]), .B(A[30]), .Y(n113) );
  NAND2XL U408 ( .A(B[8]), .B(A[8]), .Y(n222) );
  NAND2XL U409 ( .A(B[13]), .B(A[13]), .Y(n203) );
  NAND2XL U410 ( .A(B[7]), .B(A[7]), .Y(n227) );
  NAND2XL U411 ( .A(B[21]), .B(A[21]), .Y(n171) );
  NAND2XL U412 ( .A(B[36]), .B(A[36]), .Y(n63) );
  NAND2XL U413 ( .A(B[22]), .B(A[22]), .Y(n166) );
  NAND2XL U414 ( .A(n438), .B(A[38]), .Y(n45) );
  INVX2 U415 ( .A(n439), .Y(n438) );
  INVX2 U416 ( .A(B[38]), .Y(n439) );
  NOR2X1 U417 ( .A(n49), .B(n83), .Y(n47) );
  CLKINVXL U418 ( .A(n67), .Y(n69) );
  OAI21X1 U419 ( .A0(n114), .A1(n65), .B0(n66), .Y(n64) );
  NAND2XL U420 ( .A(n85), .B(n67), .Y(n65) );
  NAND2X1 U421 ( .A(n89), .B(n103), .Y(n83) );
  OAI21XL U422 ( .A0(n114), .A1(n83), .B0(n84), .Y(n82) );
  OAI21XL U423 ( .A0(n114), .A1(n101), .B0(n102), .Y(n100) );
  INVX2 U424 ( .A(n144), .Y(n143) );
  INVX2 U425 ( .A(n426), .Y(n163) );
  OAI21XL U426 ( .A0(n163), .A1(n150), .B0(n151), .Y(n149) );
  OAI21X1 U427 ( .A0(n46), .A1(n44), .B0(n45), .Y(n43) );
  NAND2XL U428 ( .A(n58), .B(n85), .Y(n56) );
  NOR2X1 U429 ( .A(n69), .B(n60), .Y(n58) );
  OAI21XL U430 ( .A0(n70), .A1(n60), .B0(n63), .Y(n59) );
  CLKINVXL U431 ( .A(n68), .Y(n70) );
  NOR2X1 U432 ( .A(n112), .B(n109), .Y(n103) );
  OAI21XL U433 ( .A0(n114), .A1(n76), .B0(n77), .Y(n75) );
  NAND2XL U434 ( .A(n85), .B(n78), .Y(n76) );
  INVX2 U435 ( .A(n81), .Y(n79) );
  NOR2X1 U436 ( .A(n125), .B(n120), .Y(n118) );
  OAI21XL U437 ( .A0(n114), .A1(n112), .B0(n113), .Y(n111) );
  NOR2X1 U438 ( .A(n141), .B(n136), .Y(n130) );
  OAI21XL U439 ( .A0(n114), .A1(n94), .B0(n95), .Y(n93) );
  NAND2XL U440 ( .A(n103), .B(n96), .Y(n94) );
  OAI21X1 U441 ( .A0(n142), .A1(n136), .B0(n137), .Y(n131) );
  NOR2X1 U442 ( .A(n150), .B(n147), .Y(n145) );
  AOI21X1 U443 ( .A0(n176), .A1(n184), .B0(n177), .Y(n175) );
  NOR2X1 U444 ( .A(n181), .B(n178), .Y(n176) );
  OAI21X1 U445 ( .A0(n178), .A1(n182), .B0(n179), .Y(n177) );
  AOI21X1 U446 ( .A0(n172), .A1(n429), .B0(n169), .Y(n167) );
  INVX2 U447 ( .A(n171), .Y(n169) );
  OAI21X1 U448 ( .A0(n173), .A1(n175), .B0(n174), .Y(n172) );
  OAI21X1 U449 ( .A0(n187), .A1(n185), .B0(n186), .Y(n184) );
  AOI21X1 U450 ( .A0(n188), .A1(n196), .B0(n189), .Y(n187) );
  OAI21X1 U451 ( .A0(n190), .A1(n194), .B0(n191), .Y(n189) );
  NOR2X1 U452 ( .A(n193), .B(n190), .Y(n188) );
  OAI21X1 U453 ( .A0(n199), .A1(n197), .B0(n198), .Y(n196) );
  AOI21X1 U454 ( .A0(n204), .A1(n430), .B0(n201), .Y(n199) );
  INVX2 U455 ( .A(n203), .Y(n201) );
  INVX2 U456 ( .A(n142), .Y(n140) );
  OAI21X1 U457 ( .A0(n221), .A1(n223), .B0(n222), .Y(n220) );
  AOI21X1 U458 ( .A0(n434), .A1(n212), .B0(n209), .Y(n207) );
  INVX2 U459 ( .A(n211), .Y(n209) );
  INVX2 U460 ( .A(n227), .Y(n225) );
  OAI21X1 U461 ( .A0(n213), .A1(n215), .B0(n214), .Y(n212) );
  AOI21X1 U462 ( .A0(n220), .A1(n436), .B0(n217), .Y(n215) );
  INVX2 U463 ( .A(n219), .Y(n217) );
  OAI21X1 U464 ( .A0(n205), .A1(n207), .B0(n206), .Y(n204) );
  AOI21X1 U465 ( .A0(n433), .A1(n240), .B0(n237), .Y(n235) );
  OAI21X1 U466 ( .A0(n229), .A1(n231), .B0(n230), .Y(n228) );
  OAI21X1 U467 ( .A0(n233), .A1(n235), .B0(n234), .Y(n232) );
  CLKINVXL U468 ( .A(n80), .Y(n78) );
  NAND2BX1 U469 ( .AN(n44), .B(n45), .Y(n2) );
  AOI21XL U470 ( .A0(n123), .A1(n143), .B0(n124), .Y(n122) );
  OAI21X1 U471 ( .A0(n133), .A1(n125), .B0(n128), .Y(n124) );
  AOI21X1 U472 ( .A0(n435), .A1(n428), .B0(n245), .Y(n243) );
  INVX2 U473 ( .A(n247), .Y(n245) );
  OAI21X1 U474 ( .A0(n241), .A1(n243), .B0(n242), .Y(n240) );
  NAND2X1 U475 ( .A(n273), .B(n431), .Y(n150) );
  NAND2BX1 U476 ( .AN(n53), .B(n54), .Y(n3) );
  NAND2BX1 U477 ( .AN(n60), .B(n63), .Y(n4) );
  OAI2BB1X1 U478 ( .A0N(n437), .A1N(n254), .B0(n253), .Y(n428) );
  NAND2XL U479 ( .A(n78), .B(n81), .Y(n6) );
  NAND2BX1 U480 ( .AN(n73), .B(n74), .Y(n5) );
  NAND2BX1 U481 ( .AN(n136), .B(n137), .Y(n13) );
  NAND2BX1 U482 ( .AN(n120), .B(n121), .Y(n11) );
  NAND2BX1 U483 ( .AN(n91), .B(n92), .Y(n7) );
  NAND2X1 U484 ( .A(n270), .B(n142), .Y(n14) );
  NAND2BX1 U485 ( .AN(n112), .B(n113), .Y(n10) );
  NAND2BX1 U486 ( .AN(n109), .B(n110), .Y(n9) );
  INVX2 U487 ( .A(n256), .Y(n254) );
  NAND2BX1 U488 ( .AN(n147), .B(n148), .Y(n15) );
  NAND2BX1 U489 ( .AN(n173), .B(n174), .Y(n20) );
  NAND2BX1 U490 ( .AN(n165), .B(n166), .Y(n18) );
  NAND2BX1 U491 ( .AN(n178), .B(n179), .Y(n21) );
  NAND2BX1 U492 ( .AN(n181), .B(n182), .Y(n22) );
  NAND2BX1 U493 ( .AN(n185), .B(n186), .Y(n23) );
  NAND2BX1 U494 ( .AN(n193), .B(n194), .Y(n25) );
  NAND2BX1 U495 ( .AN(n197), .B(n198), .Y(n26) );
  NAND2BX1 U496 ( .AN(n190), .B(n191), .Y(n24) );
  NAND2BX1 U497 ( .AN(n205), .B(n206), .Y(n28) );
  NAND2BX1 U498 ( .AN(n213), .B(n214), .Y(n30) );
  NAND2BX1 U499 ( .AN(n221), .B(n222), .Y(n32) );
  NAND2BX1 U500 ( .AN(n229), .B(n230), .Y(n34) );
  NAND2BX1 U501 ( .AN(n233), .B(n234), .Y(n35) );
  NAND2BX1 U502 ( .AN(n241), .B(n242), .Y(n37) );
  NAND2X1 U503 ( .A(n435), .B(n247), .Y(n38) );
  NAND2X1 U504 ( .A(n437), .B(n253), .Y(n39) );
  XNOR2X1 U505 ( .A(n43), .B(n1), .Y(SUM[39]) );
  XNOR2X1 U506 ( .A(n55), .B(n3), .Y(SUM[37]) );
  NOR2X1 U507 ( .A(B[37]), .B(A[37]), .Y(n53) );
  XOR2X1 U508 ( .A(n46), .B(n2), .Y(SUM[38]) );
  XNOR2X1 U509 ( .A(n64), .B(n4), .Y(SUM[36]) );
  NOR2X1 U510 ( .A(B[31]), .B(A[31]), .Y(n109) );
  NAND2XL U511 ( .A(B[35]), .B(A[35]), .Y(n74) );
  XNOR2X1 U512 ( .A(n75), .B(n5), .Y(SUM[35]) );
  NAND2XL U513 ( .A(B[37]), .B(A[37]), .Y(n54) );
  XNOR2X1 U514 ( .A(n111), .B(n9), .Y(SUM[31]) );
  NOR2X1 U515 ( .A(B[28]), .B(A[28]), .Y(n125) );
  NOR2X1 U516 ( .A(B[27]), .B(A[27]), .Y(n136) );
  XNOR2X1 U517 ( .A(n82), .B(n6), .Y(SUM[34]) );
  XNOR2X1 U518 ( .A(n100), .B(n8), .Y(SUM[32]) );
  XNOR2X1 U519 ( .A(n93), .B(n7), .Y(SUM[33]) );
  NOR2X1 U520 ( .A(B[32]), .B(A[32]), .Y(n98) );
  NOR2X1 U521 ( .A(B[30]), .B(A[30]), .Y(n112) );
  NOR2X1 U522 ( .A(B[26]), .B(A[26]), .Y(n141) );
  NOR2X1 U523 ( .A(B[15]), .B(A[15]), .Y(n193) );
  NOR2X1 U524 ( .A(B[14]), .B(A[14]), .Y(n197) );
  OR2XL U525 ( .A(B[21]), .B(A[21]), .Y(n429) );
  NOR2X1 U526 ( .A(B[20]), .B(A[20]), .Y(n173) );
  NOR2X1 U527 ( .A(B[25]), .B(A[25]), .Y(n147) );
  OR2XL U528 ( .A(B[13]), .B(A[13]), .Y(n430) );
  XOR2X1 U529 ( .A(n129), .B(n12), .Y(SUM[28]) );
  XOR2X1 U530 ( .A(n138), .B(n13), .Y(SUM[27]) );
  NOR2X1 U531 ( .A(B[19]), .B(A[19]), .Y(n178) );
  NOR2X1 U532 ( .A(B[17]), .B(A[17]), .Y(n185) );
  OR2X1 U533 ( .A(B[7]), .B(A[7]), .Y(n432) );
  NOR2X1 U534 ( .A(B[16]), .B(A[16]), .Y(n190) );
  NOR2X1 U535 ( .A(B[18]), .B(A[18]), .Y(n181) );
  NOR2X1 U536 ( .A(B[6]), .B(A[6]), .Y(n229) );
  NOR2X1 U537 ( .A(B[12]), .B(A[12]), .Y(n205) );
  NOR2X1 U538 ( .A(n438), .B(A[38]), .Y(n44) );
  NAND2XL U539 ( .A(B[14]), .B(A[14]), .Y(n198) );
  NOR2X1 U540 ( .A(B[10]), .B(A[10]), .Y(n213) );
  NOR2X1 U541 ( .A(B[5]), .B(A[5]), .Y(n233) );
  XOR2X1 U542 ( .A(n122), .B(n11), .Y(SUM[29]) );
  NAND2XL U543 ( .A(B[19]), .B(A[19]), .Y(n179) );
  OR2XL U544 ( .A(B[11]), .B(A[11]), .Y(n434) );
  NAND2XL U545 ( .A(B[24]), .B(A[24]), .Y(n155) );
  NAND2X1 U546 ( .A(B[32]), .B(A[32]), .Y(n99) );
  NAND2X1 U547 ( .A(n438), .B(A[39]), .Y(n42) );
  NOR2X1 U548 ( .A(n438), .B(A[39]), .Y(n41) );
  NAND2XL U549 ( .A(B[27]), .B(A[27]), .Y(n137) );
  NAND2XL U550 ( .A(B[20]), .B(A[20]), .Y(n174) );
  NAND2XL U551 ( .A(B[33]), .B(A[33]), .Y(n92) );
  NAND2XL U552 ( .A(B[31]), .B(A[31]), .Y(n110) );
  NAND2XL U553 ( .A(B[28]), .B(A[28]), .Y(n128) );
  OR2XL U554 ( .A(B[2]), .B(A[2]), .Y(n435) );
  NAND2XL U555 ( .A(B[25]), .B(A[25]), .Y(n148) );
  NOR2X1 U556 ( .A(B[23]), .B(A[23]), .Y(n157) );
  NAND2XL U557 ( .A(B[4]), .B(A[4]), .Y(n239) );
  OR2XL U558 ( .A(B[9]), .B(A[9]), .Y(n436) );
  NAND2XL U559 ( .A(B[29]), .B(A[29]), .Y(n121) );
  NAND2XL U560 ( .A(B[16]), .B(A[16]), .Y(n191) );
  NAND2XL U561 ( .A(B[5]), .B(A[5]), .Y(n234) );
  OR2XL U562 ( .A(B[1]), .B(A[1]), .Y(n437) );
  NAND2XL U563 ( .A(B[17]), .B(A[17]), .Y(n186) );
  NAND2XL U564 ( .A(B[11]), .B(A[11]), .Y(n211) );
  NAND2XL U565 ( .A(B[6]), .B(A[6]), .Y(n230) );
  NAND2XL U566 ( .A(B[12]), .B(A[12]), .Y(n206) );
  NAND2XL U567 ( .A(B[2]), .B(A[2]), .Y(n247) );
  NAND2XL U568 ( .A(B[10]), .B(A[10]), .Y(n214) );
  NOR2X1 U569 ( .A(B[8]), .B(A[8]), .Y(n221) );
  NOR2X1 U570 ( .A(B[3]), .B(A[3]), .Y(n241) );
  NAND2XL U571 ( .A(B[9]), .B(A[9]), .Y(n219) );
  NAND2XL U572 ( .A(B[1]), .B(A[1]), .Y(n253) );
  NAND2XL U573 ( .A(B[3]), .B(A[3]), .Y(n242) );
  XNOR2X1 U574 ( .A(n143), .B(n14), .Y(SUM[26]) );
  XNOR2X1 U575 ( .A(n156), .B(n16), .Y(SUM[24]) );
  XNOR2X1 U576 ( .A(n149), .B(n15), .Y(SUM[25]) );
  NOR2X1 U577 ( .A(B[22]), .B(A[22]), .Y(n165) );
  XOR2X1 U578 ( .A(n163), .B(n17), .Y(SUM[23]) );
  NAND2X1 U579 ( .A(B[0]), .B(A[0]), .Y(n256) );
  XOR2XL U580 ( .A(n20), .B(n175), .Y(SUM[20]) );
  XNOR2X1 U581 ( .A(n180), .B(n21), .Y(SUM[19]) );
  XOR2X1 U582 ( .A(n183), .B(n22), .Y(SUM[18]) );
  XOR2X1 U583 ( .A(n187), .B(n23), .Y(SUM[17]) );
  XNOR2X1 U584 ( .A(n192), .B(n24), .Y(SUM[16]) );
  XOR2X1 U585 ( .A(n25), .B(n195), .Y(SUM[15]) );
  XNOR2XL U586 ( .A(n27), .B(n204), .Y(SUM[13]) );
  XOR2XL U587 ( .A(n28), .B(n207), .Y(SUM[12]) );
  XNOR2XL U588 ( .A(n29), .B(n212), .Y(SUM[11]) );
  XNOR2XL U589 ( .A(n33), .B(n228), .Y(SUM[7]) );
  XOR2XL U590 ( .A(n34), .B(n231), .Y(SUM[6]) );
  XNOR2X1 U591 ( .A(n39), .B(n254), .Y(SUM[1]) );
  NAND2BX1 U592 ( .AN(n255), .B(n256), .Y(n40) );
  NOR2X1 U593 ( .A(B[0]), .B(A[0]), .Y(n255) );
  INVX2 U594 ( .A(n40), .Y(SUM[0]) );
  XOR2X1 U595 ( .A(n114), .B(n10), .Y(SUM[30]) );
  NAND2X1 U596 ( .A(n130), .B(n118), .Y(n116) );
  XNOR2X1 U597 ( .A(n172), .B(n19), .Y(SUM[21]) );
  OAI21X1 U598 ( .A0(n151), .A1(n147), .B0(n148), .Y(n146) );
  XOR2XL U599 ( .A(n32), .B(n223), .Y(SUM[8]) );
  XOR2XL U600 ( .A(n30), .B(n215), .Y(SUM[10]) );
  XOR2XL U601 ( .A(n18), .B(n167), .Y(SUM[22]) );
  XOR2XL U602 ( .A(n26), .B(n199), .Y(SUM[14]) );
endmodule


module MMSA_DW01_add_38 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n63, n64, n65, n66, n67, n68, n69, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n128, n129, n130, n131, n133, n136,
         n137, n138, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n153, n155, n156, n157, n158, n160, n163, n164,
         n165, n166, n167, n169, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n201, n203, n204, n205, n206, n207, n209, n211, n212, n213, n214,
         n215, n217, n219, n220, n221, n222, n223, n225, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n237, n239, n240, n241, n242,
         n243, n245, n247, n253, n254, n255, n256, n270, n273, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435;

  AOI21X1 U17 ( .A0(n51), .A1(n68), .B0(n52), .Y(n50) );
  AOI21X1 U27 ( .A0(n58), .A1(n86), .B0(n59), .Y(n57) );
  AOI21X1 U53 ( .A0(n86), .A1(n78), .B0(n79), .Y(n77) );
  AOI21X1 U67 ( .A0(n89), .A1(n104), .B0(n90), .Y(n84) );
  AOI21X1 U77 ( .A0(n104), .A1(n96), .B0(n97), .Y(n95) );
  AOI21X1 U108 ( .A0(n131), .A1(n118), .B0(n119), .Y(n117) );
  AOI21X1 U116 ( .A0(n123), .A1(n143), .B0(n124), .Y(n122) );
  AOI21X1 U126 ( .A0(n143), .A1(n130), .B0(n131), .Y(n129) );
  AOI21X1 U138 ( .A0(n143), .A1(n270), .B0(n140), .Y(n138) );
  AOI21X1 U157 ( .A0(n427), .A1(n160), .B0(n153), .Y(n151) );
  AOI21X1 U217 ( .A0(n188), .A1(n196), .B0(n189), .Y(n187) );
  AOI21X1 U252 ( .A0(n431), .A1(n212), .B0(n209), .Y(n207) );
  AOI21X1 U266 ( .A0(n220), .A1(n425), .B0(n217), .Y(n215) );
  AOI21X1 U315 ( .A0(n432), .A1(n424), .B0(n245), .Y(n243) );
  NOR2XL U340 ( .A(B[34]), .B(A[34]), .Y(n80) );
  XNOR2X2 U341 ( .A(n43), .B(n1), .Y(SUM[39]) );
  OAI21X2 U342 ( .A0(n46), .A1(n44), .B0(n45), .Y(n43) );
  NOR2XL U343 ( .A(n49), .B(n83), .Y(n47) );
  NOR2XL U344 ( .A(B[35]), .B(A[35]), .Y(n73) );
  CLKINVXL U345 ( .A(n84), .Y(n86) );
  AOI21XL U346 ( .A0(n86), .A1(n67), .B0(n68), .Y(n66) );
  INVX1 U347 ( .A(n67), .Y(n69) );
  AOI21X1 U348 ( .A0(n145), .A1(n164), .B0(n146), .Y(n144) );
  NOR2X1 U349 ( .A(n91), .B(n98), .Y(n89) );
  NOR2X1 U350 ( .A(B[19]), .B(A[19]), .Y(n178) );
  OAI21X1 U351 ( .A0(n109), .A1(n113), .B0(n110), .Y(n104) );
  OAI21X1 U352 ( .A0(n73), .A1(n81), .B0(n74), .Y(n68) );
  NOR2X1 U353 ( .A(n60), .B(n53), .Y(n51) );
  NOR2X1 U354 ( .A(n80), .B(n73), .Y(n67) );
  OAI21X2 U355 ( .A0(n116), .A1(n144), .B0(n117), .Y(n115) );
  NOR2X1 U356 ( .A(n125), .B(n120), .Y(n118) );
  NOR2X1 U357 ( .A(B[25]), .B(A[25]), .Y(n147) );
  NOR2X1 U358 ( .A(B[28]), .B(A[28]), .Y(n125) );
  NOR2X1 U359 ( .A(B[31]), .B(A[31]), .Y(n109) );
  NOR2X1 U360 ( .A(B[29]), .B(A[29]), .Y(n120) );
  NOR2X1 U361 ( .A(B[36]), .B(A[36]), .Y(n60) );
  OAI21XL U362 ( .A0(n114), .A1(n83), .B0(n84), .Y(n82) );
  OAI21X2 U363 ( .A0(n165), .A1(n167), .B0(n166), .Y(n164) );
  OAI21X1 U364 ( .A0(n84), .A1(n49), .B0(n50), .Y(n48) );
  INVX1 U365 ( .A(n155), .Y(n153) );
  OAI21XL U366 ( .A0(n53), .A1(n63), .B0(n54), .Y(n52) );
  CLKINVX2 U367 ( .A(n158), .Y(n160) );
  NAND2BXL U368 ( .AN(n109), .B(n110), .Y(n9) );
  NAND2BX1 U369 ( .AN(n41), .B(n42), .Y(n1) );
  NOR2X1 U370 ( .A(B[27]), .B(A[27]), .Y(n136) );
  OAI21XL U371 ( .A0(n114), .A1(n101), .B0(n102), .Y(n100) );
  CLKINVXL U372 ( .A(n103), .Y(n101) );
  NAND2XL U373 ( .A(n103), .B(n96), .Y(n94) );
  OAI21XL U374 ( .A0(n114), .A1(n56), .B0(n57), .Y(n55) );
  OAI21XL U375 ( .A0(n114), .A1(n76), .B0(n77), .Y(n75) );
  CLKINVXL U376 ( .A(n81), .Y(n79) );
  CLKINVXL U377 ( .A(n60), .Y(n423) );
  NAND2BX1 U378 ( .AN(n91), .B(n92), .Y(n7) );
  CLKINVX2 U379 ( .A(n211), .Y(n209) );
  NAND2BX1 U380 ( .AN(n73), .B(n74), .Y(n5) );
  NAND2X1 U381 ( .A(B[30]), .B(A[30]), .Y(n113) );
  OR2XL U382 ( .A(B[9]), .B(A[9]), .Y(n425) );
  NAND2XL U383 ( .A(n89), .B(n103), .Y(n83) );
  CLKINVXL U384 ( .A(n144), .Y(n143) );
  INVX1 U385 ( .A(n115), .Y(n114) );
  CLKINVXL U386 ( .A(n164), .Y(n163) );
  OAI21XL U387 ( .A0(n163), .A1(n150), .B0(n151), .Y(n149) );
  CLKINVXL U388 ( .A(n131), .Y(n133) );
  CLKINVXL U389 ( .A(n184), .Y(n183) );
  AOI21X1 U390 ( .A0(n172), .A1(n426), .B0(n169), .Y(n167) );
  NOR2BXL U391 ( .AN(n130), .B(n125), .Y(n123) );
  CLKINVXL U392 ( .A(n99), .Y(n97) );
  OAI21X1 U393 ( .A0(n199), .A1(n197), .B0(n198), .Y(n196) );
  CLKINVX1 U394 ( .A(n219), .Y(n217) );
  CLKINVXL U395 ( .A(n98), .Y(n96) );
  OAI21X1 U396 ( .A0(n120), .A1(n128), .B0(n121), .Y(n119) );
  NOR2X1 U397 ( .A(n112), .B(n109), .Y(n103) );
  CLKINVX2 U398 ( .A(n157), .Y(n273) );
  NAND2XL U399 ( .A(n96), .B(n99), .Y(n8) );
  OAI2BB1X1 U400 ( .A0N(n68), .A1N(n423), .B0(n63), .Y(n59) );
  INVX1 U401 ( .A(n232), .Y(n231) );
  NAND2XL U402 ( .A(n427), .B(n155), .Y(n16) );
  CLKINVXL U403 ( .A(n141), .Y(n270) );
  CLKINVXL U404 ( .A(n80), .Y(n78) );
  NAND2BXL U405 ( .AN(n125), .B(n128), .Y(n12) );
  NAND2BXL U406 ( .AN(n178), .B(n179), .Y(n21) );
  OAI21XL U407 ( .A0(n183), .A1(n181), .B0(n182), .Y(n180) );
  NAND2BXL U408 ( .AN(n181), .B(n182), .Y(n22) );
  OAI21XL U409 ( .A0(n195), .A1(n193), .B0(n194), .Y(n192) );
  NAND2XL U410 ( .A(n431), .B(n211), .Y(n29) );
  OR2XL U411 ( .A(B[24]), .B(A[24]), .Y(n427) );
  NAND2XL U412 ( .A(B[27]), .B(A[27]), .Y(n137) );
  NAND2XL U413 ( .A(B[26]), .B(A[26]), .Y(n142) );
  NAND2XL U414 ( .A(B[15]), .B(A[15]), .Y(n194) );
  NAND2XL U415 ( .A(B[8]), .B(A[8]), .Y(n222) );
  OR2XL U416 ( .A(B[13]), .B(A[13]), .Y(n429) );
  NAND2XL U417 ( .A(B[20]), .B(A[20]), .Y(n174) );
  NOR2X1 U418 ( .A(B[33]), .B(A[33]), .Y(n91) );
  NAND2XL U419 ( .A(B[13]), .B(A[13]), .Y(n203) );
  OR2XL U420 ( .A(B[7]), .B(A[7]), .Y(n430) );
  OR2XL U421 ( .A(B[21]), .B(A[21]), .Y(n426) );
  NAND2XL U422 ( .A(B[23]), .B(A[23]), .Y(n158) );
  NAND2XL U423 ( .A(B[21]), .B(A[21]), .Y(n171) );
  NAND2XL U424 ( .A(B[14]), .B(A[14]), .Y(n198) );
  NAND2XL U425 ( .A(B[7]), .B(A[7]), .Y(n227) );
  NAND2XL U426 ( .A(B[34]), .B(A[34]), .Y(n81) );
  NAND2XL U427 ( .A(B[36]), .B(A[36]), .Y(n63) );
  NAND2XL U428 ( .A(B[22]), .B(A[22]), .Y(n166) );
  NAND2XL U429 ( .A(n434), .B(A[38]), .Y(n45) );
  INVX2 U430 ( .A(n435), .Y(n434) );
  INVX2 U431 ( .A(B[38]), .Y(n435) );
  INVX2 U432 ( .A(n83), .Y(n85) );
  AOI21X1 U433 ( .A0(n115), .A1(n47), .B0(n48), .Y(n46) );
  NAND2X1 U434 ( .A(n67), .B(n51), .Y(n49) );
  OAI21XL U435 ( .A0(n114), .A1(n65), .B0(n66), .Y(n64) );
  CLKINVXL U436 ( .A(n104), .Y(n102) );
  INVX2 U437 ( .A(n196), .Y(n195) );
  NAND2XL U438 ( .A(n58), .B(n85), .Y(n56) );
  NOR2X1 U439 ( .A(n69), .B(n60), .Y(n58) );
  NAND2X1 U440 ( .A(n130), .B(n118), .Y(n116) );
  OAI21X1 U441 ( .A0(n91), .A1(n99), .B0(n92), .Y(n90) );
  AOI21X1 U442 ( .A0(n176), .A1(n184), .B0(n177), .Y(n175) );
  OAI21X1 U443 ( .A0(n178), .A1(n182), .B0(n179), .Y(n177) );
  NOR2X1 U444 ( .A(n181), .B(n178), .Y(n176) );
  OAI21X1 U445 ( .A0(n151), .A1(n147), .B0(n148), .Y(n146) );
  NOR2X1 U446 ( .A(n150), .B(n147), .Y(n145) );
  OAI21X1 U447 ( .A0(n173), .A1(n175), .B0(n174), .Y(n172) );
  INVX2 U448 ( .A(n171), .Y(n169) );
  OAI21X1 U449 ( .A0(n142), .A1(n136), .B0(n137), .Y(n131) );
  OAI21X1 U450 ( .A0(n190), .A1(n194), .B0(n191), .Y(n189) );
  NOR2X1 U451 ( .A(n193), .B(n190), .Y(n188) );
  AOI21X1 U452 ( .A0(n204), .A1(n429), .B0(n201), .Y(n199) );
  INVX2 U453 ( .A(n203), .Y(n201) );
  OAI21X1 U454 ( .A0(n205), .A1(n207), .B0(n206), .Y(n204) );
  OAI21X1 U455 ( .A0(n213), .A1(n215), .B0(n214), .Y(n212) );
  OAI21X1 U456 ( .A0(n187), .A1(n185), .B0(n186), .Y(n184) );
  NAND2XL U457 ( .A(n85), .B(n78), .Y(n76) );
  NOR2X1 U458 ( .A(n141), .B(n136), .Y(n130) );
  OAI21XL U459 ( .A0(n114), .A1(n112), .B0(n113), .Y(n111) );
  OAI21XL U460 ( .A0(n133), .A1(n125), .B0(n128), .Y(n124) );
  OAI21XL U461 ( .A0(n114), .A1(n94), .B0(n95), .Y(n93) );
  INVX2 U462 ( .A(n142), .Y(n140) );
  AOI21X1 U463 ( .A0(n228), .A1(n430), .B0(n225), .Y(n223) );
  INVX2 U464 ( .A(n227), .Y(n225) );
  OAI21X1 U465 ( .A0(n229), .A1(n231), .B0(n230), .Y(n228) );
  OAI21X1 U466 ( .A0(n221), .A1(n223), .B0(n222), .Y(n220) );
  OAI21X1 U467 ( .A0(n233), .A1(n235), .B0(n234), .Y(n232) );
  AOI21X1 U468 ( .A0(n428), .A1(n240), .B0(n237), .Y(n235) );
  NAND2X1 U469 ( .A(n273), .B(n427), .Y(n150) );
  NAND2BX1 U470 ( .AN(n44), .B(n45), .Y(n2) );
  OAI21X1 U471 ( .A0(n241), .A1(n243), .B0(n242), .Y(n240) );
  INVX2 U472 ( .A(n247), .Y(n245) );
  NAND2BX1 U473 ( .AN(n53), .B(n54), .Y(n3) );
  NAND2BX1 U474 ( .AN(n60), .B(n63), .Y(n4) );
  OAI2BB1X1 U475 ( .A0N(n433), .A1N(n254), .B0(n253), .Y(n424) );
  NAND2XL U476 ( .A(n78), .B(n81), .Y(n6) );
  OAI21X1 U477 ( .A0(n163), .A1(n157), .B0(n158), .Y(n156) );
  NAND2BX1 U478 ( .AN(n120), .B(n121), .Y(n11) );
  NAND2BX1 U479 ( .AN(n112), .B(n113), .Y(n10) );
  NAND2X1 U480 ( .A(n270), .B(n142), .Y(n14) );
  NAND2BX1 U481 ( .AN(n147), .B(n148), .Y(n15) );
  NAND2BX1 U482 ( .AN(n136), .B(n137), .Y(n13) );
  INVX2 U483 ( .A(n256), .Y(n254) );
  NAND2XL U484 ( .A(n273), .B(n158), .Y(n17) );
  NAND2BX1 U485 ( .AN(n173), .B(n174), .Y(n20) );
  NAND2X1 U486 ( .A(n426), .B(n171), .Y(n19) );
  NAND2BX1 U487 ( .AN(n165), .B(n166), .Y(n18) );
  NAND2BX1 U488 ( .AN(n185), .B(n186), .Y(n23) );
  NAND2BX1 U489 ( .AN(n190), .B(n191), .Y(n24) );
  NAND2BX1 U490 ( .AN(n193), .B(n194), .Y(n25) );
  NAND2BX1 U491 ( .AN(n197), .B(n198), .Y(n26) );
  NAND2X1 U492 ( .A(n429), .B(n203), .Y(n27) );
  NAND2BX1 U493 ( .AN(n205), .B(n206), .Y(n28) );
  NAND2BX1 U494 ( .AN(n213), .B(n214), .Y(n30) );
  NAND2XL U495 ( .A(n425), .B(n219), .Y(n31) );
  NAND2BX1 U496 ( .AN(n221), .B(n222), .Y(n32) );
  NAND2X1 U497 ( .A(n430), .B(n227), .Y(n33) );
  NAND2BX1 U498 ( .AN(n229), .B(n230), .Y(n34) );
  NAND2BX1 U499 ( .AN(n233), .B(n234), .Y(n35) );
  NAND2BX1 U500 ( .AN(n241), .B(n242), .Y(n37) );
  NAND2X1 U501 ( .A(n432), .B(n247), .Y(n38) );
  NAND2X1 U502 ( .A(n433), .B(n253), .Y(n39) );
  NOR2X1 U503 ( .A(B[37]), .B(A[37]), .Y(n53) );
  XNOR2X1 U504 ( .A(n55), .B(n3), .Y(SUM[37]) );
  NAND2XL U505 ( .A(B[35]), .B(A[35]), .Y(n74) );
  NAND2XL U506 ( .A(B[37]), .B(A[37]), .Y(n54) );
  XNOR2X1 U507 ( .A(n82), .B(n6), .Y(SUM[34]) );
  NOR2X1 U508 ( .A(B[20]), .B(A[20]), .Y(n173) );
  NOR2X1 U509 ( .A(B[18]), .B(A[18]), .Y(n181) );
  NOR2X1 U510 ( .A(B[16]), .B(A[16]), .Y(n190) );
  XNOR2X1 U511 ( .A(n64), .B(n4), .Y(SUM[36]) );
  XNOR2X1 U512 ( .A(n75), .B(n5), .Y(SUM[35]) );
  NOR2X1 U513 ( .A(B[14]), .B(A[14]), .Y(n197) );
  NOR2X1 U514 ( .A(B[26]), .B(A[26]), .Y(n141) );
  XNOR2X1 U515 ( .A(n111), .B(n9), .Y(SUM[31]) );
  XOR2X1 U516 ( .A(n122), .B(n11), .Y(SUM[29]) );
  XNOR2X1 U517 ( .A(n93), .B(n7), .Y(SUM[33]) );
  NAND2X1 U518 ( .A(B[18]), .B(A[18]), .Y(n182) );
  XNOR2X1 U519 ( .A(n100), .B(n8), .Y(SUM[32]) );
  XOR2X1 U520 ( .A(n129), .B(n12), .Y(SUM[28]) );
  XOR2X1 U521 ( .A(n138), .B(n13), .Y(SUM[27]) );
  NOR2X1 U522 ( .A(B[15]), .B(A[15]), .Y(n193) );
  NOR2X1 U523 ( .A(B[12]), .B(A[12]), .Y(n205) );
  NOR2X1 U524 ( .A(B[32]), .B(A[32]), .Y(n98) );
  NOR2X1 U525 ( .A(B[5]), .B(A[5]), .Y(n233) );
  OR2XL U526 ( .A(B[4]), .B(A[4]), .Y(n428) );
  XOR2X1 U527 ( .A(n114), .B(n10), .Y(SUM[30]) );
  NOR2X1 U528 ( .A(B[17]), .B(A[17]), .Y(n185) );
  NAND2XL U529 ( .A(B[28]), .B(A[28]), .Y(n128) );
  NAND2XL U530 ( .A(B[19]), .B(A[19]), .Y(n179) );
  NOR2X1 U531 ( .A(B[6]), .B(A[6]), .Y(n229) );
  NOR2X1 U532 ( .A(B[23]), .B(A[23]), .Y(n157) );
  NOR2X1 U533 ( .A(n434), .B(A[38]), .Y(n44) );
  NAND2X1 U534 ( .A(B[32]), .B(A[32]), .Y(n99) );
  OR2XL U535 ( .A(B[11]), .B(A[11]), .Y(n431) );
  NAND2XL U536 ( .A(B[29]), .B(A[29]), .Y(n121) );
  NOR2X1 U537 ( .A(B[30]), .B(A[30]), .Y(n112) );
  NOR2X1 U538 ( .A(B[10]), .B(A[10]), .Y(n213) );
  NAND2XL U539 ( .A(B[16]), .B(A[16]), .Y(n191) );
  NAND2XL U540 ( .A(B[31]), .B(A[31]), .Y(n110) );
  NAND2XL U541 ( .A(B[24]), .B(A[24]), .Y(n155) );
  NAND2XL U542 ( .A(B[12]), .B(A[12]), .Y(n206) );
  NAND2XL U543 ( .A(B[5]), .B(A[5]), .Y(n234) );
  NAND2XL U544 ( .A(B[33]), .B(A[33]), .Y(n92) );
  NAND2XL U545 ( .A(B[25]), .B(A[25]), .Y(n148) );
  NAND2XL U546 ( .A(B[11]), .B(A[11]), .Y(n211) );
  OR2XL U547 ( .A(B[2]), .B(A[2]), .Y(n432) );
  NAND2XL U548 ( .A(B[17]), .B(A[17]), .Y(n186) );
  NAND2X1 U549 ( .A(n434), .B(A[39]), .Y(n42) );
  NOR2X1 U550 ( .A(n434), .B(A[39]), .Y(n41) );
  NOR2X1 U551 ( .A(B[3]), .B(A[3]), .Y(n241) );
  NOR2X1 U552 ( .A(B[8]), .B(A[8]), .Y(n221) );
  NAND2XL U553 ( .A(B[6]), .B(A[6]), .Y(n230) );
  NAND2XL U554 ( .A(B[2]), .B(A[2]), .Y(n247) );
  NAND2XL U555 ( .A(B[10]), .B(A[10]), .Y(n214) );
  OR2XL U556 ( .A(B[1]), .B(A[1]), .Y(n433) );
  XNOR2X1 U557 ( .A(n143), .B(n14), .Y(SUM[26]) );
  NAND2XL U558 ( .A(B[3]), .B(A[3]), .Y(n242) );
  NAND2XL U559 ( .A(B[1]), .B(A[1]), .Y(n253) );
  NOR2X1 U560 ( .A(B[22]), .B(A[22]), .Y(n165) );
  XNOR2X1 U561 ( .A(n149), .B(n15), .Y(SUM[25]) );
  XNOR2X1 U562 ( .A(n156), .B(n16), .Y(SUM[24]) );
  XOR2X1 U563 ( .A(n163), .B(n17), .Y(SUM[23]) );
  NAND2X1 U564 ( .A(B[0]), .B(A[0]), .Y(n256) );
  XNOR2X1 U565 ( .A(n172), .B(n19), .Y(SUM[21]) );
  XNOR2X1 U566 ( .A(n180), .B(n21), .Y(SUM[19]) );
  XOR2X1 U567 ( .A(n183), .B(n22), .Y(SUM[18]) );
  XNOR2X1 U568 ( .A(n192), .B(n24), .Y(SUM[16]) );
  XOR2X1 U569 ( .A(n25), .B(n195), .Y(SUM[15]) );
  XOR2XL U570 ( .A(n26), .B(n199), .Y(SUM[14]) );
  XNOR2XL U571 ( .A(n29), .B(n212), .Y(SUM[11]) );
  XNOR2XL U572 ( .A(n31), .B(n220), .Y(SUM[9]) );
  XOR2XL U573 ( .A(n32), .B(n223), .Y(SUM[8]) );
  XNOR2XL U574 ( .A(n33), .B(n228), .Y(SUM[7]) );
  XOR2XL U575 ( .A(n34), .B(n231), .Y(SUM[6]) );
  XOR2XL U576 ( .A(n35), .B(n235), .Y(SUM[5]) );
  XNOR2X1 U577 ( .A(n38), .B(n424), .Y(SUM[2]) );
  XNOR2X1 U578 ( .A(n39), .B(n254), .Y(SUM[1]) );
  NAND2BX1 U579 ( .AN(n255), .B(n256), .Y(n40) );
  NOR2X1 U580 ( .A(B[0]), .B(A[0]), .Y(n255) );
  INVX2 U581 ( .A(n40), .Y(SUM[0]) );
  NAND2XL U582 ( .A(n428), .B(n239), .Y(n36) );
  CLKINVX2 U583 ( .A(n239), .Y(n237) );
  NAND2XL U584 ( .A(B[4]), .B(A[4]), .Y(n239) );
  NAND2XL U585 ( .A(n85), .B(n67), .Y(n65) );
  XNOR2XL U586 ( .A(n27), .B(n204), .Y(SUM[13]) );
  XOR2X1 U587 ( .A(n187), .B(n23), .Y(SUM[17]) );
  NAND2XL U588 ( .A(B[9]), .B(A[9]), .Y(n219) );
  XOR2XL U589 ( .A(n18), .B(n167), .Y(SUM[22]) );
  XOR2XL U590 ( .A(n20), .B(n175), .Y(SUM[20]) );
  XNOR2XL U591 ( .A(n36), .B(n240), .Y(SUM[4]) );
  XOR2XL U592 ( .A(n37), .B(n243), .Y(SUM[3]) );
  XOR2XL U593 ( .A(n28), .B(n207), .Y(SUM[12]) );
  XOR2XL U594 ( .A(n30), .B(n215), .Y(SUM[10]) );
  XOR2X1 U595 ( .A(n46), .B(n2), .Y(SUM[38]) );
endmodule


module MMSA_DW01_add_37 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n20, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n63,
         n64, n65, n66, n67, n68, n70, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n128, n129, n130, n131, n133, n136, n137, n138, n140,
         n141, n142, n144, n145, n146, n147, n148, n149, n150, n151, n153,
         n155, n156, n157, n158, n160, n163, n164, n165, n166, n167, n169,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n201, n203, n204, n205,
         n206, n207, n209, n211, n212, n213, n214, n215, n217, n219, n220,
         n221, n222, n223, n225, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n237, n239, n240, n241, n242, n243, n245, n247, n253,
         n254, n255, n256, n258, n259, n260, n263, n267, n268, n270, n271,
         n273, n276, n277, n278, n281, n282, n286, n290, n293, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441;

  AOI21X1 U17 ( .A0(n51), .A1(n68), .B0(n52), .Y(n50) );
  AOI21X1 U27 ( .A0(n58), .A1(n86), .B0(n59), .Y(n57) );
  AOI21X1 U39 ( .A0(n86), .A1(n67), .B0(n68), .Y(n66) );
  AOI21X1 U53 ( .A0(n86), .A1(n78), .B0(n79), .Y(n77) );
  AOI21X1 U77 ( .A0(n104), .A1(n96), .B0(n97), .Y(n95) );
  AOI21X1 U126 ( .A0(n424), .A1(n130), .B0(n131), .Y(n129) );
  AOI21X1 U138 ( .A0(n424), .A1(n270), .B0(n140), .Y(n138) );
  AOI21X1 U157 ( .A0(n435), .A1(n160), .B0(n153), .Y(n151) );
  AOI21X1 U266 ( .A0(n220), .A1(n438), .B0(n217), .Y(n215) );
  AOI21X1 U301 ( .A0(n431), .A1(n240), .B0(n237), .Y(n235) );
  AOI21X1 U315 ( .A0(n432), .A1(n430), .B0(n245), .Y(n243) );
  CLKINVX2 U340 ( .A(n116), .Y(n423) );
  NAND2X1 U341 ( .A(n130), .B(n118), .Y(n116) );
  NOR2X1 U342 ( .A(n125), .B(n120), .Y(n118) );
  NOR2X1 U343 ( .A(B[6]), .B(A[6]), .Y(n229) );
  NOR2X1 U344 ( .A(B[19]), .B(A[19]), .Y(n178) );
  NOR2X1 U345 ( .A(B[18]), .B(A[18]), .Y(n181) );
  NOR2X1 U346 ( .A(n60), .B(n53), .Y(n51) );
  NAND2X2 U347 ( .A(n425), .B(n117), .Y(n115) );
  AOI21X1 U348 ( .A0(n131), .A1(n118), .B0(n119), .Y(n117) );
  NAND2X1 U349 ( .A(n423), .B(n424), .Y(n425) );
  NOR2X1 U350 ( .A(n80), .B(n73), .Y(n67) );
  NOR2X1 U351 ( .A(B[36]), .B(A[36]), .Y(n60) );
  INVX2 U352 ( .A(n115), .Y(n114) );
  AOI21X1 U353 ( .A0(n145), .A1(n164), .B0(n146), .Y(n144) );
  CLKINVX2 U354 ( .A(n144), .Y(n424) );
  OAI21X1 U355 ( .A0(n114), .A1(n101), .B0(n102), .Y(n100) );
  AOI21XL U356 ( .A0(n115), .A1(n47), .B0(n48), .Y(n46) );
  NOR2BX1 U357 ( .AN(n67), .B(n60), .Y(n58) );
  OAI21XL U358 ( .A0(n73), .A1(n81), .B0(n74), .Y(n68) );
  CLKINVX1 U359 ( .A(n155), .Y(n153) );
  NAND2XL U360 ( .A(n58), .B(n85), .Y(n56) );
  OAI21XL U361 ( .A0(n53), .A1(n63), .B0(n54), .Y(n52) );
  OAI21XL U362 ( .A0(n114), .A1(n65), .B0(n66), .Y(n64) );
  NAND2XL U363 ( .A(n78), .B(n81), .Y(n6) );
  CLKINVX1 U364 ( .A(n158), .Y(n160) );
  NAND2BX1 U365 ( .AN(n136), .B(n137), .Y(n13) );
  INVX1 U366 ( .A(n44), .Y(n258) );
  CLKINVXL U367 ( .A(n241), .Y(n293) );
  OAI21XL U368 ( .A0(n84), .A1(n49), .B0(n50), .Y(n48) );
  NAND2XL U369 ( .A(n89), .B(n103), .Y(n83) );
  CLKINVXL U370 ( .A(n104), .Y(n102) );
  CLKINVXL U371 ( .A(n103), .Y(n101) );
  CLKINVXL U372 ( .A(n131), .Y(n133) );
  OAI21XL U373 ( .A0(n163), .A1(n150), .B0(n151), .Y(n149) );
  CLKINVXL U374 ( .A(n184), .Y(n183) );
  CLKINVXL U375 ( .A(n196), .Y(n195) );
  OAI21X1 U376 ( .A0(n70), .A1(n60), .B0(n63), .Y(n59) );
  NAND2XL U377 ( .A(n260), .B(n63), .Y(n4) );
  OAI21XL U378 ( .A0(n151), .A1(n147), .B0(n148), .Y(n146) );
  CLKINVXL U379 ( .A(n99), .Y(n97) );
  NAND2XL U380 ( .A(n103), .B(n96), .Y(n94) );
  NAND2XL U381 ( .A(n263), .B(n92), .Y(n7) );
  XOR2X1 U382 ( .A(n100), .B(n426), .Y(SUM[32]) );
  AND2X1 U383 ( .A(n96), .B(n99), .Y(n426) );
  AOI21X1 U384 ( .A0(n172), .A1(n434), .B0(n169), .Y(n167) );
  NOR2BXL U385 ( .AN(n130), .B(n125), .Y(n123) );
  NAND2XL U386 ( .A(n267), .B(n121), .Y(n11) );
  NAND2XL U387 ( .A(n268), .B(n128), .Y(n12) );
  CLKINVXL U388 ( .A(n98), .Y(n96) );
  CLKINVX1 U389 ( .A(n219), .Y(n217) );
  OAI21XL U390 ( .A0(n163), .A1(n157), .B0(n158), .Y(n156) );
  XOR2X1 U391 ( .A(n156), .B(n427), .Y(SUM[24]) );
  AND2X1 U392 ( .A(n435), .B(n155), .Y(n427) );
  NAND2XL U393 ( .A(n271), .B(n148), .Y(n15) );
  CLKINVX2 U394 ( .A(n157), .Y(n273) );
  INVX1 U395 ( .A(n232), .Y(n231) );
  CLKINVXL U396 ( .A(n141), .Y(n270) );
  CLKINVXL U397 ( .A(n147), .Y(n271) );
  CLKINVXL U398 ( .A(n91), .Y(n263) );
  XOR2X1 U399 ( .A(n172), .B(n428), .Y(SUM[21]) );
  AND2X1 U400 ( .A(n434), .B(n171), .Y(n428) );
  CLKINVXL U401 ( .A(n80), .Y(n78) );
  CLKINVXL U402 ( .A(n53), .Y(n259) );
  NAND2XL U403 ( .A(n276), .B(n174), .Y(n20) );
  CLKINVXL U404 ( .A(n173), .Y(n276) );
  XOR2X1 U405 ( .A(n180), .B(n429), .Y(SUM[19]) );
  AND2X1 U406 ( .A(n277), .B(n179), .Y(n429) );
  OAI21XL U407 ( .A0(n195), .A1(n193), .B0(n194), .Y(n192) );
  CLKINVXL U408 ( .A(n193), .Y(n281) );
  NAND2XL U409 ( .A(n282), .B(n198), .Y(n26) );
  CLKINVXL U410 ( .A(n197), .Y(n282) );
  NAND2XL U411 ( .A(n437), .B(n203), .Y(n27) );
  NAND2XL U412 ( .A(n439), .B(n211), .Y(n29) );
  NAND2XL U413 ( .A(n286), .B(n214), .Y(n30) );
  CLKINVXL U414 ( .A(n213), .Y(n286) );
  NAND2XL U415 ( .A(n438), .B(n219), .Y(n31) );
  OR2XL U416 ( .A(B[24]), .B(A[24]), .Y(n435) );
  NOR2X1 U417 ( .A(B[27]), .B(A[27]), .Y(n136) );
  NAND2XL U418 ( .A(B[26]), .B(A[26]), .Y(n142) );
  NAND2XL U419 ( .A(B[18]), .B(A[18]), .Y(n182) );
  NAND2XL U420 ( .A(B[15]), .B(A[15]), .Y(n194) );
  NAND2XL U421 ( .A(B[8]), .B(A[8]), .Y(n222) );
  NAND2XL U422 ( .A(B[30]), .B(A[30]), .Y(n113) );
  OR2XL U423 ( .A(B[21]), .B(A[21]), .Y(n434) );
  OR2XL U424 ( .A(B[7]), .B(A[7]), .Y(n433) );
  NAND2XL U425 ( .A(B[23]), .B(A[23]), .Y(n158) );
  NAND2XL U426 ( .A(B[7]), .B(A[7]), .Y(n227) );
  NAND2XL U427 ( .A(B[21]), .B(A[21]), .Y(n171) );
  NAND2XL U428 ( .A(B[6]), .B(A[6]), .Y(n230) );
  NOR2X1 U429 ( .A(B[30]), .B(A[30]), .Y(n112) );
  NOR2X1 U430 ( .A(B[29]), .B(A[29]), .Y(n120) );
  NAND2XL U431 ( .A(B[34]), .B(A[34]), .Y(n81) );
  NAND2XL U432 ( .A(B[22]), .B(A[22]), .Y(n166) );
  OR2XL U433 ( .A(B[4]), .B(A[4]), .Y(n431) );
  NAND2XL U434 ( .A(B[4]), .B(A[4]), .Y(n239) );
  NAND2BX1 U435 ( .AN(n41), .B(n42), .Y(n1) );
  NAND2XL U436 ( .A(n440), .B(A[38]), .Y(n45) );
  INVX2 U437 ( .A(n441), .Y(n440) );
  INVX2 U438 ( .A(B[38]), .Y(n441) );
  INVX2 U439 ( .A(n83), .Y(n85) );
  NOR2X1 U440 ( .A(n49), .B(n83), .Y(n47) );
  NAND2X1 U441 ( .A(n67), .B(n51), .Y(n49) );
  INVX2 U442 ( .A(n68), .Y(n70) );
  NAND2X1 U443 ( .A(n85), .B(n67), .Y(n65) );
  OAI21XL U444 ( .A0(n114), .A1(n83), .B0(n84), .Y(n82) );
  INVX2 U445 ( .A(n164), .Y(n163) );
  OAI21X1 U446 ( .A0(n46), .A1(n44), .B0(n45), .Y(n43) );
  NAND2X1 U447 ( .A(n259), .B(n54), .Y(n3) );
  XOR2X1 U448 ( .A(n46), .B(n2), .Y(SUM[38]) );
  NAND2X1 U449 ( .A(n258), .B(n45), .Y(n2) );
  AOI21X1 U450 ( .A0(n228), .A1(n433), .B0(n225), .Y(n223) );
  INVX2 U451 ( .A(n227), .Y(n225) );
  OAI21X1 U452 ( .A0(n241), .A1(n243), .B0(n242), .Y(n240) );
  AOI21X1 U453 ( .A0(n439), .A1(n212), .B0(n209), .Y(n207) );
  INVX2 U454 ( .A(n211), .Y(n209) );
  AOI21X1 U455 ( .A0(n176), .A1(n184), .B0(n177), .Y(n175) );
  OAI21X1 U456 ( .A0(n178), .A1(n182), .B0(n179), .Y(n177) );
  NOR2X1 U457 ( .A(n181), .B(n178), .Y(n176) );
  INVX2 U458 ( .A(n239), .Y(n237) );
  OAI21X1 U459 ( .A0(n213), .A1(n215), .B0(n214), .Y(n212) );
  CLKINVX2 U460 ( .A(n247), .Y(n245) );
  AOI21X1 U461 ( .A0(n204), .A1(n437), .B0(n201), .Y(n199) );
  INVX2 U462 ( .A(n203), .Y(n201) );
  OAI21X1 U463 ( .A0(n187), .A1(n185), .B0(n186), .Y(n184) );
  OAI21X1 U464 ( .A0(n165), .A1(n167), .B0(n166), .Y(n164) );
  OAI21X1 U465 ( .A0(n199), .A1(n197), .B0(n198), .Y(n196) );
  OAI21X1 U466 ( .A0(n205), .A1(n207), .B0(n206), .Y(n204) );
  OAI21X1 U467 ( .A0(n229), .A1(n231), .B0(n230), .Y(n228) );
  AOI21X1 U468 ( .A0(n188), .A1(n196), .B0(n189), .Y(n187) );
  OAI21X1 U469 ( .A0(n190), .A1(n194), .B0(n191), .Y(n189) );
  NOR2X1 U470 ( .A(n193), .B(n190), .Y(n188) );
  OAI21X1 U471 ( .A0(n173), .A1(n175), .B0(n174), .Y(n172) );
  OAI21X1 U472 ( .A0(n221), .A1(n223), .B0(n222), .Y(n220) );
  NOR2X1 U473 ( .A(n150), .B(n147), .Y(n145) );
  INVX2 U474 ( .A(n171), .Y(n169) );
  OAI21X1 U475 ( .A0(n233), .A1(n235), .B0(n234), .Y(n232) );
  XOR2X1 U476 ( .A(n129), .B(n12), .Y(SUM[28]) );
  OAI21X1 U477 ( .A0(n142), .A1(n136), .B0(n137), .Y(n131) );
  XNOR2X1 U478 ( .A(n64), .B(n4), .Y(SUM[36]) );
  AOI21XL U479 ( .A0(n123), .A1(n424), .B0(n124), .Y(n122) );
  XOR2X1 U480 ( .A(n122), .B(n11), .Y(SUM[29]) );
  INVX2 U481 ( .A(n142), .Y(n140) );
  OAI21XL U482 ( .A0(n114), .A1(n94), .B0(n95), .Y(n93) );
  XNOR2X1 U483 ( .A(n93), .B(n7), .Y(SUM[33]) );
  NOR2X1 U484 ( .A(n141), .B(n136), .Y(n130) );
  NOR2X1 U485 ( .A(n112), .B(n109), .Y(n103) );
  NOR2X1 U486 ( .A(n91), .B(n98), .Y(n89) );
  OAI21XL U487 ( .A0(n114), .A1(n76), .B0(n77), .Y(n75) );
  NAND2XL U488 ( .A(n85), .B(n78), .Y(n76) );
  INVX2 U489 ( .A(n81), .Y(n79) );
  XNOR2X1 U490 ( .A(n82), .B(n6), .Y(SUM[34]) );
  OAI21XL U491 ( .A0(n114), .A1(n112), .B0(n113), .Y(n111) );
  OAI21X1 U492 ( .A0(n120), .A1(n128), .B0(n121), .Y(n119) );
  OAI2BB1X1 U493 ( .A0N(n436), .A1N(n254), .B0(n253), .Y(n430) );
  AOI21X1 U494 ( .A0(n89), .A1(n104), .B0(n90), .Y(n84) );
  NAND2X1 U495 ( .A(n273), .B(n435), .Y(n150) );
  OAI21X1 U496 ( .A0(n109), .A1(n113), .B0(n110), .Y(n104) );
  CLKINVXL U497 ( .A(n60), .Y(n260) );
  XNOR2X1 U498 ( .A(n149), .B(n15), .Y(SUM[25]) );
  NAND2BX1 U499 ( .AN(n73), .B(n74), .Y(n5) );
  INVX2 U500 ( .A(n256), .Y(n254) );
  NAND2X1 U501 ( .A(n270), .B(n142), .Y(n14) );
  INVX2 U502 ( .A(n120), .Y(n267) );
  NAND2BX1 U503 ( .AN(n112), .B(n113), .Y(n10) );
  NAND2BX1 U504 ( .AN(n109), .B(n110), .Y(n9) );
  XOR2XL U505 ( .A(n20), .B(n175), .Y(SUM[20]) );
  NAND2XL U506 ( .A(n273), .B(n158), .Y(n17) );
  NAND2BX1 U507 ( .AN(n165), .B(n166), .Y(n18) );
  OAI21XL U508 ( .A0(n183), .A1(n181), .B0(n182), .Y(n180) );
  XOR2X1 U509 ( .A(n183), .B(n22), .Y(SUM[18]) );
  NAND2X1 U510 ( .A(n278), .B(n182), .Y(n22) );
  CLKINVXL U511 ( .A(n181), .Y(n278) );
  CLKINVXL U512 ( .A(n178), .Y(n277) );
  NAND2BX1 U513 ( .AN(n185), .B(n186), .Y(n23) );
  XOR2X1 U514 ( .A(n25), .B(n195), .Y(SUM[15]) );
  NAND2X1 U515 ( .A(n281), .B(n194), .Y(n25) );
  NAND2BX1 U516 ( .AN(n190), .B(n191), .Y(n24) );
  NAND2BX1 U517 ( .AN(n205), .B(n206), .Y(n28) );
  XNOR2XL U518 ( .A(n29), .B(n212), .Y(SUM[11]) );
  NAND2BX1 U519 ( .AN(n221), .B(n222), .Y(n32) );
  XNOR2XL U520 ( .A(n33), .B(n228), .Y(SUM[7]) );
  NAND2X1 U521 ( .A(n433), .B(n227), .Y(n33) );
  CLKINVXL U522 ( .A(n229), .Y(n290) );
  XOR2XL U523 ( .A(n34), .B(n231), .Y(SUM[6]) );
  NAND2X1 U524 ( .A(n290), .B(n230), .Y(n34) );
  NAND2BX1 U525 ( .AN(n233), .B(n234), .Y(n35) );
  NAND2X1 U526 ( .A(n431), .B(n239), .Y(n36) );
  NAND2X1 U527 ( .A(n293), .B(n242), .Y(n37) );
  XNOR2XL U528 ( .A(n38), .B(n430), .Y(SUM[2]) );
  NAND2XL U529 ( .A(n432), .B(n247), .Y(n38) );
  NAND2X1 U530 ( .A(n436), .B(n253), .Y(n39) );
  NOR2X1 U531 ( .A(B[37]), .B(A[37]), .Y(n53) );
  XNOR2X1 U532 ( .A(n43), .B(n1), .Y(SUM[39]) );
  NOR2X1 U533 ( .A(B[35]), .B(A[35]), .Y(n73) );
  NOR2X1 U534 ( .A(B[34]), .B(A[34]), .Y(n80) );
  NOR2X1 U535 ( .A(B[28]), .B(A[28]), .Y(n125) );
  NAND2XL U536 ( .A(B[36]), .B(A[36]), .Y(n63) );
  NOR2X1 U537 ( .A(B[14]), .B(A[14]), .Y(n197) );
  NAND2XL U538 ( .A(B[35]), .B(A[35]), .Y(n74) );
  NAND2XL U539 ( .A(B[37]), .B(A[37]), .Y(n54) );
  NOR2X1 U540 ( .A(B[5]), .B(A[5]), .Y(n233) );
  NOR2X1 U541 ( .A(B[20]), .B(A[20]), .Y(n173) );
  XOR2X1 U542 ( .A(n138), .B(n13), .Y(SUM[27]) );
  OR2X1 U543 ( .A(B[2]), .B(A[2]), .Y(n432) );
  NOR2X1 U544 ( .A(B[31]), .B(A[31]), .Y(n109) );
  NOR2X1 U545 ( .A(B[25]), .B(A[25]), .Y(n147) );
  NOR2X1 U546 ( .A(B[26]), .B(A[26]), .Y(n141) );
  NOR2X1 U547 ( .A(B[32]), .B(A[32]), .Y(n98) );
  NOR2X1 U548 ( .A(B[15]), .B(A[15]), .Y(n193) );
  NAND2XL U549 ( .A(B[27]), .B(A[27]), .Y(n137) );
  NOR2X1 U550 ( .A(B[16]), .B(A[16]), .Y(n190) );
  NOR2X1 U551 ( .A(B[3]), .B(A[3]), .Y(n241) );
  XNOR2X1 U552 ( .A(n75), .B(n5), .Y(SUM[35]) );
  XNOR2X1 U553 ( .A(n111), .B(n9), .Y(SUM[31]) );
  NOR2X1 U554 ( .A(B[17]), .B(A[17]), .Y(n185) );
  NOR2X1 U555 ( .A(B[12]), .B(A[12]), .Y(n205) );
  NAND2XL U556 ( .A(B[14]), .B(A[14]), .Y(n198) );
  NOR2X1 U557 ( .A(B[33]), .B(A[33]), .Y(n91) );
  OR2X1 U558 ( .A(B[1]), .B(A[1]), .Y(n436) );
  NAND2XL U559 ( .A(B[28]), .B(A[28]), .Y(n128) );
  NAND2XL U560 ( .A(B[20]), .B(A[20]), .Y(n174) );
  NAND2X1 U561 ( .A(B[32]), .B(A[32]), .Y(n99) );
  NAND2XL U562 ( .A(B[5]), .B(A[5]), .Y(n234) );
  OR2XL U563 ( .A(B[13]), .B(A[13]), .Y(n437) );
  NAND2XL U564 ( .A(B[19]), .B(A[19]), .Y(n179) );
  XOR2X1 U565 ( .A(n114), .B(n10), .Y(SUM[30]) );
  NAND2XL U566 ( .A(B[29]), .B(A[29]), .Y(n121) );
  NOR2X1 U567 ( .A(B[23]), .B(A[23]), .Y(n157) );
  OR2XL U568 ( .A(B[9]), .B(A[9]), .Y(n438) );
  NAND2XL U569 ( .A(B[16]), .B(A[16]), .Y(n191) );
  NOR2X1 U570 ( .A(B[10]), .B(A[10]), .Y(n213) );
  NAND2XL U571 ( .A(B[24]), .B(A[24]), .Y(n155) );
  OR2XL U572 ( .A(B[11]), .B(A[11]), .Y(n439) );
  NAND2XL U573 ( .A(B[13]), .B(A[13]), .Y(n203) );
  NAND2X1 U574 ( .A(B[1]), .B(A[1]), .Y(n253) );
  NAND2XL U575 ( .A(B[33]), .B(A[33]), .Y(n92) );
  NAND2XL U576 ( .A(B[12]), .B(A[12]), .Y(n206) );
  NAND2XL U577 ( .A(B[17]), .B(A[17]), .Y(n186) );
  NAND2XL U578 ( .A(B[3]), .B(A[3]), .Y(n242) );
  NAND2XL U579 ( .A(B[25]), .B(A[25]), .Y(n148) );
  NOR2X1 U580 ( .A(n440), .B(A[38]), .Y(n44) );
  NAND2XL U581 ( .A(B[11]), .B(A[11]), .Y(n211) );
  NAND2XL U582 ( .A(B[9]), .B(A[9]), .Y(n219) );
  NOR2X1 U583 ( .A(B[8]), .B(A[8]), .Y(n221) );
  NAND2XL U584 ( .A(B[31]), .B(A[31]), .Y(n110) );
  NAND2X1 U585 ( .A(n440), .B(A[39]), .Y(n42) );
  NOR2X1 U586 ( .A(n440), .B(A[39]), .Y(n41) );
  NAND2XL U587 ( .A(B[10]), .B(A[10]), .Y(n214) );
  XNOR2X1 U588 ( .A(n424), .B(n14), .Y(SUM[26]) );
  NOR2X1 U589 ( .A(B[22]), .B(A[22]), .Y(n165) );
  XOR2X1 U590 ( .A(n163), .B(n17), .Y(SUM[23]) );
  NAND2X1 U591 ( .A(B[0]), .B(A[0]), .Y(n256) );
  XOR2X1 U592 ( .A(n187), .B(n23), .Y(SUM[17]) );
  XNOR2X1 U593 ( .A(n192), .B(n24), .Y(SUM[16]) );
  XNOR2XL U594 ( .A(n27), .B(n204), .Y(SUM[13]) );
  XOR2XL U595 ( .A(n28), .B(n207), .Y(SUM[12]) );
  XNOR2XL U596 ( .A(n31), .B(n220), .Y(SUM[9]) );
  XOR2XL U597 ( .A(n32), .B(n223), .Y(SUM[8]) );
  XNOR2XL U598 ( .A(n36), .B(n240), .Y(SUM[4]) );
  XNOR2X1 U599 ( .A(n39), .B(n254), .Y(SUM[1]) );
  NAND2BX1 U600 ( .AN(n255), .B(n256), .Y(n40) );
  NOR2X1 U601 ( .A(B[0]), .B(A[0]), .Y(n255) );
  INVX2 U602 ( .A(n40), .Y(SUM[0]) );
  OAI21XL U603 ( .A0(n133), .A1(n125), .B0(n128), .Y(n124) );
  CLKINVXL U604 ( .A(n125), .Y(n268) );
  XNOR2X1 U605 ( .A(n55), .B(n3), .Y(SUM[37]) );
  OAI21X1 U606 ( .A0(n91), .A1(n99), .B0(n92), .Y(n90) );
  OAI21X1 U607 ( .A0(n114), .A1(n56), .B0(n57), .Y(n55) );
  INVX2 U608 ( .A(n84), .Y(n86) );
  XOR2XL U609 ( .A(n30), .B(n215), .Y(SUM[10]) );
  XOR2XL U610 ( .A(n18), .B(n167), .Y(SUM[22]) );
  XOR2XL U611 ( .A(n37), .B(n243), .Y(SUM[3]) );
  XOR2XL U612 ( .A(n26), .B(n199), .Y(SUM[14]) );
  XOR2XL U613 ( .A(n35), .B(n235), .Y(SUM[5]) );
  NAND2X1 U614 ( .A(B[2]), .B(A[2]), .Y(n247) );
endmodule


module MMSA_DW01_add_36 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n63, n64, n66, n67, n68, n69, n70, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n128, n129, n130, n131, n132, n133, n136, n137,
         n138, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n153, n155, n156, n157, n158, n160, n163, n164, n165,
         n166, n167, n169, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n201,
         n203, n204, n205, n206, n207, n209, n211, n212, n213, n214, n215,
         n217, n219, n220, n221, n222, n223, n225, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n237, n239, n240, n241, n242, n243,
         n245, n247, n253, n254, n255, n256, n258, n259, n260, n263, n267,
         n268, n270, n271, n273, n276, n277, n278, n281, n282, n286, n290,
         n293, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436;

  AOI21X1 U13 ( .A0(n115), .A1(n47), .B0(n48), .Y(n46) );
  AOI21X1 U17 ( .A0(n51), .A1(n68), .B0(n52), .Y(n50) );
  AOI21X1 U27 ( .A0(n58), .A1(n86), .B0(n59), .Y(n57) );
  AOI21X1 U39 ( .A0(n86), .A1(n67), .B0(n68), .Y(n66) );
  AOI21X1 U53 ( .A0(n86), .A1(n78), .B0(n79), .Y(n77) );
  AOI21X1 U77 ( .A0(n104), .A1(n96), .B0(n97), .Y(n95) );
  AOI21X1 U108 ( .A0(n131), .A1(n118), .B0(n119), .Y(n117) );
  AOI21X1 U138 ( .A0(n143), .A1(n270), .B0(n140), .Y(n138) );
  AOI21X1 U157 ( .A0(n431), .A1(n160), .B0(n153), .Y(n151) );
  AOI21X1 U217 ( .A0(n188), .A1(n196), .B0(n189), .Y(n187) );
  AOI21X1 U266 ( .A0(n220), .A1(n435), .B0(n217), .Y(n215) );
  AOI21X1 U280 ( .A0(n228), .A1(n434), .B0(n225), .Y(n223) );
  AOI21X1 U315 ( .A0(n433), .A1(n427), .B0(n245), .Y(n243) );
  AOI21X1 U340 ( .A0(n145), .A1(n164), .B0(n146), .Y(n144) );
  OAI21X1 U341 ( .A0(n116), .A1(n144), .B0(n117), .Y(n115) );
  NAND2X1 U342 ( .A(n130), .B(n118), .Y(n116) );
  NOR2X1 U343 ( .A(n112), .B(n109), .Y(n103) );
  NOR2X1 U344 ( .A(B[29]), .B(A[29]), .Y(n120) );
  NOR2X1 U345 ( .A(B[27]), .B(A[27]), .Y(n136) );
  NOR2X1 U346 ( .A(B[30]), .B(A[30]), .Y(n112) );
  NOR2X1 U347 ( .A(n49), .B(n83), .Y(n47) );
  OAI2BB1X1 U348 ( .A0N(n115), .A1N(n423), .B0(n66), .Y(n64) );
  AND2X1 U349 ( .A(n85), .B(n67), .Y(n423) );
  INVX2 U350 ( .A(n115), .Y(n114) );
  INVXL U351 ( .A(n155), .Y(n153) );
  INVXL U352 ( .A(n67), .Y(n69) );
  AOI21XL U353 ( .A0(n143), .A1(n130), .B0(n131), .Y(n129) );
  INVXL U354 ( .A(n68), .Y(n70) );
  NAND2XL U355 ( .A(n89), .B(n103), .Y(n83) );
  OAI21X1 U356 ( .A0(n114), .A1(n56), .B0(n57), .Y(n55) );
  NAND2X1 U357 ( .A(n58), .B(n85), .Y(n56) );
  OAI21XL U358 ( .A0(n53), .A1(n63), .B0(n54), .Y(n52) );
  NOR2X1 U359 ( .A(B[33]), .B(A[33]), .Y(n91) );
  OR2XL U360 ( .A(B[24]), .B(A[24]), .Y(n431) );
  INVXL U361 ( .A(n103), .Y(n101) );
  OAI21XL U362 ( .A0(n114), .A1(n76), .B0(n77), .Y(n75) );
  CLKINVXL U363 ( .A(n81), .Y(n79) );
  CLKINVX1 U364 ( .A(n158), .Y(n160) );
  INVX1 U365 ( .A(n44), .Y(n258) );
  NAND2BX1 U366 ( .AN(n73), .B(n74), .Y(n5) );
  NAND2XL U367 ( .A(n429), .B(n171), .Y(n19) );
  CLKINVXL U368 ( .A(n241), .Y(n293) );
  OAI21XL U369 ( .A0(n84), .A1(n49), .B0(n50), .Y(n48) );
  CLKINVXL U370 ( .A(n104), .Y(n102) );
  CLKINVXL U371 ( .A(n164), .Y(n163) );
  OAI21XL U372 ( .A0(n163), .A1(n150), .B0(n151), .Y(n149) );
  CLKINVXL U373 ( .A(n130), .Y(n132) );
  CLKINVXL U374 ( .A(n184), .Y(n183) );
  CLKINVXL U375 ( .A(n196), .Y(n195) );
  CLKINVXL U376 ( .A(n99), .Y(n97) );
  OAI21X1 U377 ( .A0(n120), .A1(n128), .B0(n121), .Y(n119) );
  NAND2XL U378 ( .A(n263), .B(n92), .Y(n7) );
  XOR2X1 U379 ( .A(n100), .B(n424), .Y(SUM[32]) );
  AND2X1 U380 ( .A(n96), .B(n99), .Y(n424) );
  NAND2XL U381 ( .A(n268), .B(n128), .Y(n12) );
  OAI21XL U382 ( .A0(n133), .A1(n125), .B0(n128), .Y(n124) );
  NAND2XL U383 ( .A(n267), .B(n121), .Y(n11) );
  NAND2XL U384 ( .A(n78), .B(n81), .Y(n6) );
  CLKINVXL U385 ( .A(n98), .Y(n96) );
  OAI21XL U386 ( .A0(n163), .A1(n157), .B0(n158), .Y(n156) );
  XOR2X1 U387 ( .A(n156), .B(n425), .Y(SUM[24]) );
  AND2X1 U388 ( .A(n431), .B(n155), .Y(n425) );
  NAND2XL U389 ( .A(n271), .B(n148), .Y(n15) );
  CLKINVX1 U390 ( .A(n219), .Y(n217) );
  CLKINVX1 U391 ( .A(n227), .Y(n225) );
  CLKINVX2 U392 ( .A(n157), .Y(n273) );
  INVX1 U393 ( .A(n232), .Y(n231) );
  CLKINVXL U394 ( .A(n141), .Y(n270) );
  CLKINVXL U395 ( .A(n147), .Y(n271) );
  CLKINVXL U396 ( .A(n125), .Y(n268) );
  CLKINVXL U397 ( .A(n60), .Y(n260) );
  CLKINVXL U398 ( .A(n53), .Y(n259) );
  NAND2XL U399 ( .A(n276), .B(n174), .Y(n20) );
  NAND2XL U400 ( .A(n273), .B(n158), .Y(n17) );
  CLKINVXL U401 ( .A(n173), .Y(n276) );
  XOR2X1 U402 ( .A(n180), .B(n426), .Y(SUM[19]) );
  AND2X1 U403 ( .A(n277), .B(n179), .Y(n426) );
  CLKINVXL U404 ( .A(n178), .Y(n277) );
  OAI21XL U405 ( .A0(n183), .A1(n181), .B0(n182), .Y(n180) );
  CLKINVXL U406 ( .A(n181), .Y(n278) );
  OAI21XL U407 ( .A0(n195), .A1(n193), .B0(n194), .Y(n192) );
  CLKINVXL U408 ( .A(n193), .Y(n281) );
  NAND2XL U409 ( .A(n282), .B(n198), .Y(n26) );
  CLKINVXL U410 ( .A(n197), .Y(n282) );
  NAND2XL U411 ( .A(n430), .B(n203), .Y(n27) );
  NAND2XL U412 ( .A(n436), .B(n211), .Y(n29) );
  NAND2XL U413 ( .A(n286), .B(n214), .Y(n30) );
  CLKINVXL U414 ( .A(n213), .Y(n286) );
  NAND2XL U415 ( .A(n435), .B(n219), .Y(n31) );
  NAND2XL U416 ( .A(n434), .B(n227), .Y(n33) );
  NAND2XL U417 ( .A(n290), .B(n230), .Y(n34) );
  CLKINVXL U418 ( .A(n229), .Y(n290) );
  NAND2XL U419 ( .A(B[26]), .B(A[26]), .Y(n142) );
  NAND2XL U420 ( .A(B[18]), .B(A[18]), .Y(n182) );
  NAND2XL U421 ( .A(B[30]), .B(A[30]), .Y(n113) );
  NAND2XL U422 ( .A(B[15]), .B(A[15]), .Y(n194) );
  NAND2XL U423 ( .A(B[8]), .B(A[8]), .Y(n222) );
  NAND2XL U424 ( .A(B[23]), .B(A[23]), .Y(n158) );
  OR2XL U425 ( .A(B[13]), .B(A[13]), .Y(n430) );
  NOR2XL U426 ( .A(B[35]), .B(A[35]), .Y(n73) );
  OR2XL U427 ( .A(B[21]), .B(A[21]), .Y(n429) );
  NAND2XL U428 ( .A(B[21]), .B(A[21]), .Y(n171) );
  NAND2XL U429 ( .A(B[34]), .B(A[34]), .Y(n81) );
  NOR2XL U430 ( .A(B[34]), .B(A[34]), .Y(n80) );
  NAND2XL U431 ( .A(B[36]), .B(A[36]), .Y(n63) );
  NAND2XL U432 ( .A(B[22]), .B(A[22]), .Y(n166) );
  NAND2BX1 U433 ( .AN(n41), .B(n42), .Y(n1) );
  INVX2 U434 ( .A(n83), .Y(n85) );
  NAND2X1 U435 ( .A(n67), .B(n51), .Y(n49) );
  OAI21XL U436 ( .A0(n114), .A1(n101), .B0(n102), .Y(n100) );
  OAI21XL U437 ( .A0(n114), .A1(n83), .B0(n84), .Y(n82) );
  INVX2 U438 ( .A(n84), .Y(n86) );
  NOR2X1 U439 ( .A(n80), .B(n73), .Y(n67) );
  NOR2X1 U440 ( .A(n69), .B(n60), .Y(n58) );
  XNOR2X1 U441 ( .A(n55), .B(n3), .Y(SUM[37]) );
  NAND2X1 U442 ( .A(n259), .B(n54), .Y(n3) );
  NOR2X1 U443 ( .A(n60), .B(n53), .Y(n51) );
  OAI21X1 U444 ( .A0(n73), .A1(n81), .B0(n74), .Y(n68) );
  NAND2X1 U445 ( .A(n258), .B(n45), .Y(n2) );
  XNOR2X1 U446 ( .A(n64), .B(n4), .Y(SUM[36]) );
  NAND2X1 U447 ( .A(n260), .B(n63), .Y(n4) );
  OAI21X1 U448 ( .A0(n70), .A1(n60), .B0(n63), .Y(n59) );
  NOR2X1 U449 ( .A(n141), .B(n136), .Y(n130) );
  OAI21XL U450 ( .A0(n114), .A1(n94), .B0(n95), .Y(n93) );
  NAND2XL U451 ( .A(n103), .B(n96), .Y(n94) );
  XNOR2X1 U452 ( .A(n93), .B(n7), .Y(SUM[33]) );
  OAI21X1 U453 ( .A0(n142), .A1(n136), .B0(n137), .Y(n131) );
  NOR2X1 U454 ( .A(n125), .B(n120), .Y(n118) );
  OAI21XL U455 ( .A0(n114), .A1(n112), .B0(n113), .Y(n111) );
  NAND2XL U456 ( .A(n85), .B(n78), .Y(n76) );
  XNOR2X1 U457 ( .A(n82), .B(n6), .Y(SUM[34]) );
  OAI21X1 U458 ( .A0(n190), .A1(n194), .B0(n191), .Y(n189) );
  NOR2X1 U459 ( .A(n193), .B(n190), .Y(n188) );
  OAI21X1 U460 ( .A0(n187), .A1(n185), .B0(n186), .Y(n184) );
  OAI21X1 U461 ( .A0(n173), .A1(n175), .B0(n174), .Y(n172) );
  AOI21X1 U462 ( .A0(n172), .A1(n429), .B0(n169), .Y(n167) );
  INVX2 U463 ( .A(n171), .Y(n169) );
  OAI21X1 U464 ( .A0(n199), .A1(n197), .B0(n198), .Y(n196) );
  OAI21X1 U465 ( .A0(n165), .A1(n167), .B0(n166), .Y(n164) );
  OAI21X1 U466 ( .A0(n151), .A1(n147), .B0(n148), .Y(n146) );
  NOR2X1 U467 ( .A(n150), .B(n147), .Y(n145) );
  AOI21X1 U468 ( .A0(n176), .A1(n184), .B0(n177), .Y(n175) );
  OAI21X1 U469 ( .A0(n178), .A1(n182), .B0(n179), .Y(n177) );
  NOR2X1 U470 ( .A(n181), .B(n178), .Y(n176) );
  AOI21X1 U471 ( .A0(n89), .A1(n104), .B0(n90), .Y(n84) );
  OAI21X1 U472 ( .A0(n91), .A1(n99), .B0(n92), .Y(n90) );
  OAI21X1 U473 ( .A0(n109), .A1(n113), .B0(n110), .Y(n104) );
  AOI21X1 U474 ( .A0(n204), .A1(n430), .B0(n201), .Y(n199) );
  INVX2 U475 ( .A(n203), .Y(n201) );
  OAI21X1 U476 ( .A0(n205), .A1(n207), .B0(n206), .Y(n204) );
  OAI21X1 U477 ( .A0(n213), .A1(n215), .B0(n214), .Y(n212) );
  OAI21X1 U478 ( .A0(n221), .A1(n223), .B0(n222), .Y(n220) );
  OAI21X1 U479 ( .A0(n229), .A1(n231), .B0(n230), .Y(n228) );
  AOI21X1 U480 ( .A0(n428), .A1(n240), .B0(n237), .Y(n235) );
  INVX2 U481 ( .A(n239), .Y(n237) );
  AOI21X1 U482 ( .A0(n436), .A1(n212), .B0(n209), .Y(n207) );
  INVX2 U483 ( .A(n211), .Y(n209) );
  OAI21X1 U484 ( .A0(n233), .A1(n235), .B0(n234), .Y(n232) );
  AOI21X1 U485 ( .A0(n123), .A1(n143), .B0(n124), .Y(n122) );
  NOR2X1 U486 ( .A(n132), .B(n125), .Y(n123) );
  CLKINVXL U487 ( .A(n131), .Y(n133) );
  XOR2X1 U488 ( .A(n129), .B(n12), .Y(SUM[28]) );
  NOR2X1 U489 ( .A(n91), .B(n98), .Y(n89) );
  INVX2 U490 ( .A(n142), .Y(n140) );
  INVX2 U491 ( .A(n247), .Y(n245) );
  OAI21X1 U492 ( .A0(n241), .A1(n243), .B0(n242), .Y(n240) );
  OAI2BB1X1 U493 ( .A0N(n432), .A1N(n254), .B0(n253), .Y(n427) );
  INVX2 U494 ( .A(n80), .Y(n78) );
  NAND2X1 U495 ( .A(n273), .B(n431), .Y(n150) );
  XNOR2X1 U496 ( .A(n149), .B(n15), .Y(SUM[25]) );
  CLKINVXL U497 ( .A(n120), .Y(n267) );
  NAND2BX1 U498 ( .AN(n136), .B(n137), .Y(n13) );
  INVX2 U499 ( .A(n256), .Y(n254) );
  INVX2 U500 ( .A(n91), .Y(n263) );
  NAND2BX1 U501 ( .AN(n112), .B(n113), .Y(n10) );
  NAND2BX1 U502 ( .AN(n109), .B(n110), .Y(n9) );
  NAND2X1 U503 ( .A(n270), .B(n142), .Y(n14) );
  XOR2X1 U504 ( .A(n183), .B(n22), .Y(SUM[18]) );
  NAND2X1 U505 ( .A(n278), .B(n182), .Y(n22) );
  NAND2BX1 U506 ( .AN(n165), .B(n166), .Y(n18) );
  NAND2BX1 U507 ( .AN(n185), .B(n186), .Y(n23) );
  XOR2X1 U508 ( .A(n25), .B(n195), .Y(SUM[15]) );
  NAND2X1 U509 ( .A(n281), .B(n194), .Y(n25) );
  XOR2XL U510 ( .A(n26), .B(n199), .Y(SUM[14]) );
  NAND2BX1 U511 ( .AN(n190), .B(n191), .Y(n24) );
  NAND2BX1 U512 ( .AN(n205), .B(n206), .Y(n28) );
  NAND2BX1 U513 ( .AN(n221), .B(n222), .Y(n32) );
  XNOR2XL U514 ( .A(n33), .B(n228), .Y(SUM[7]) );
  XOR2XL U515 ( .A(n34), .B(n231), .Y(SUM[6]) );
  NAND2XL U516 ( .A(n428), .B(n239), .Y(n36) );
  NAND2BX1 U517 ( .AN(n233), .B(n234), .Y(n35) );
  XOR2X1 U518 ( .A(n37), .B(n243), .Y(SUM[3]) );
  NAND2X1 U519 ( .A(n293), .B(n242), .Y(n37) );
  XNOR2X1 U520 ( .A(n38), .B(n427), .Y(SUM[2]) );
  NAND2X1 U521 ( .A(n432), .B(n253), .Y(n39) );
  XNOR2X1 U522 ( .A(n43), .B(n1), .Y(SUM[39]) );
  NOR2X1 U523 ( .A(B[37]), .B(A[37]), .Y(n53) );
  NOR2X1 U524 ( .A(B[36]), .B(A[36]), .Y(n60) );
  NAND2XL U525 ( .A(B[35]), .B(A[35]), .Y(n74) );
  NAND2XL U526 ( .A(B[37]), .B(A[37]), .Y(n54) );
  NOR2X1 U527 ( .A(B[31]), .B(A[31]), .Y(n109) );
  NOR2X1 U528 ( .A(B[28]), .B(A[28]), .Y(n125) );
  XNOR2X1 U529 ( .A(n111), .B(n9), .Y(SUM[31]) );
  XNOR2X1 U530 ( .A(n75), .B(n5), .Y(SUM[35]) );
  NOR2X1 U531 ( .A(B[14]), .B(A[14]), .Y(n197) );
  NOR2X1 U532 ( .A(B[26]), .B(A[26]), .Y(n141) );
  NOR2X1 U533 ( .A(B[19]), .B(A[19]), .Y(n178) );
  NOR2X1 U534 ( .A(B[18]), .B(A[18]), .Y(n181) );
  NOR2X1 U535 ( .A(B[20]), .B(A[20]), .Y(n173) );
  OR2XL U536 ( .A(B[4]), .B(A[4]), .Y(n428) );
  XOR2X1 U537 ( .A(n114), .B(n10), .Y(SUM[30]) );
  NOR2X1 U538 ( .A(B[32]), .B(A[32]), .Y(n98) );
  NOR2X1 U539 ( .A(B[16]), .B(A[16]), .Y(n190) );
  NOR2X1 U540 ( .A(B[15]), .B(A[15]), .Y(n193) );
  NOR2X1 U541 ( .A(B[25]), .B(A[25]), .Y(n147) );
  NAND2XL U542 ( .A(B[14]), .B(A[14]), .Y(n198) );
  NAND2XL U543 ( .A(B[27]), .B(A[27]), .Y(n137) );
  NOR2X1 U544 ( .A(B[38]), .B(A[38]), .Y(n44) );
  NOR2X1 U545 ( .A(B[17]), .B(A[17]), .Y(n185) );
  NOR2X1 U546 ( .A(B[12]), .B(A[12]), .Y(n205) );
  NAND2XL U547 ( .A(B[28]), .B(A[28]), .Y(n128) );
  NAND2XL U548 ( .A(B[20]), .B(A[20]), .Y(n174) );
  NAND2X1 U549 ( .A(B[32]), .B(A[32]), .Y(n99) );
  NOR2X1 U550 ( .A(B[5]), .B(A[5]), .Y(n233) );
  NAND2XL U551 ( .A(B[31]), .B(A[31]), .Y(n110) );
  NAND2XL U552 ( .A(B[33]), .B(A[33]), .Y(n92) );
  NAND2XL U553 ( .A(B[19]), .B(A[19]), .Y(n179) );
  OR2XL U554 ( .A(B[1]), .B(A[1]), .Y(n432) );
  OR2XL U555 ( .A(B[2]), .B(A[2]), .Y(n433) );
  NAND2XL U556 ( .A(B[16]), .B(A[16]), .Y(n191) );
  NAND2XL U557 ( .A(B[13]), .B(A[13]), .Y(n203) );
  NAND2XL U558 ( .A(B[29]), .B(A[29]), .Y(n121) );
  OR2XL U559 ( .A(B[7]), .B(A[7]), .Y(n434) );
  NAND2XL U560 ( .A(B[12]), .B(A[12]), .Y(n206) );
  NOR2X1 U561 ( .A(B[6]), .B(A[6]), .Y(n229) );
  NAND2XL U562 ( .A(B[38]), .B(A[39]), .Y(n42) );
  NOR2X1 U563 ( .A(B[38]), .B(A[39]), .Y(n41) );
  NOR2X1 U564 ( .A(B[23]), .B(A[23]), .Y(n157) );
  NOR2X1 U565 ( .A(B[10]), .B(A[10]), .Y(n213) );
  NAND2XL U566 ( .A(B[38]), .B(A[38]), .Y(n45) );
  NAND2XL U567 ( .A(B[24]), .B(A[24]), .Y(n155) );
  OR2XL U568 ( .A(B[9]), .B(A[9]), .Y(n435) );
  NAND2XL U569 ( .A(B[11]), .B(A[11]), .Y(n211) );
  OR2XL U570 ( .A(B[11]), .B(A[11]), .Y(n436) );
  NAND2XL U571 ( .A(B[17]), .B(A[17]), .Y(n186) );
  NAND2XL U572 ( .A(B[5]), .B(A[5]), .Y(n234) );
  NAND2XL U573 ( .A(B[1]), .B(A[1]), .Y(n253) );
  NAND2XL U574 ( .A(B[7]), .B(A[7]), .Y(n227) );
  NAND2XL U575 ( .A(B[25]), .B(A[25]), .Y(n148) );
  XNOR2X1 U576 ( .A(n143), .B(n14), .Y(SUM[26]) );
  NAND2XL U577 ( .A(B[9]), .B(A[9]), .Y(n219) );
  NAND2XL U578 ( .A(B[6]), .B(A[6]), .Y(n230) );
  NOR2X1 U579 ( .A(B[8]), .B(A[8]), .Y(n221) );
  NAND2XL U580 ( .A(B[10]), .B(A[10]), .Y(n214) );
  NOR2X1 U581 ( .A(B[3]), .B(A[3]), .Y(n241) );
  XOR2X1 U582 ( .A(n163), .B(n17), .Y(SUM[23]) );
  NOR2X1 U583 ( .A(B[22]), .B(A[22]), .Y(n165) );
  NAND2XL U584 ( .A(B[3]), .B(A[3]), .Y(n242) );
  NAND2X1 U585 ( .A(B[0]), .B(A[0]), .Y(n256) );
  XOR2XL U586 ( .A(n18), .B(n167), .Y(SUM[22]) );
  XNOR2X1 U587 ( .A(n192), .B(n24), .Y(SUM[16]) );
  XNOR2XL U588 ( .A(n31), .B(n220), .Y(SUM[9]) );
  XNOR2X1 U589 ( .A(n39), .B(n254), .Y(SUM[1]) );
  NAND2BX1 U590 ( .AN(n255), .B(n256), .Y(n40) );
  NOR2X1 U591 ( .A(B[0]), .B(A[0]), .Y(n255) );
  INVX2 U592 ( .A(n40), .Y(SUM[0]) );
  NAND2XL U593 ( .A(B[4]), .B(A[4]), .Y(n239) );
  XNOR2XL U594 ( .A(n29), .B(n212), .Y(SUM[11]) );
  XOR2XL U595 ( .A(n35), .B(n235), .Y(SUM[5]) );
  XNOR2XL U596 ( .A(n27), .B(n204), .Y(SUM[13]) );
  XNOR2X1 U597 ( .A(n172), .B(n19), .Y(SUM[21]) );
  XOR2X1 U598 ( .A(n138), .B(n13), .Y(SUM[27]) );
  XOR2X1 U599 ( .A(n122), .B(n11), .Y(SUM[29]) );
  XOR2XL U600 ( .A(n20), .B(n175), .Y(SUM[20]) );
  INVX2 U601 ( .A(n144), .Y(n143) );
  XOR2XL U602 ( .A(n28), .B(n207), .Y(SUM[12]) );
  XOR2X1 U603 ( .A(n46), .B(n2), .Y(SUM[38]) );
  XOR2XL U604 ( .A(n30), .B(n215), .Y(SUM[10]) );
  XNOR2XL U605 ( .A(n36), .B(n240), .Y(SUM[4]) );
  NAND2XL U606 ( .A(n433), .B(n247), .Y(n38) );
  XOR2X1 U607 ( .A(n187), .B(n23), .Y(SUM[17]) );
  XOR2XL U608 ( .A(n32), .B(n223), .Y(SUM[8]) );
  OAI21X1 U609 ( .A0(n46), .A1(n44), .B0(n45), .Y(n43) );
  NAND2X1 U610 ( .A(B[2]), .B(A[2]), .Y(n247) );
endmodule


module MMSA_DW01_add_35 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n63,
         n64, n65, n66, n67, n68, n70, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n128, n129, n130, n131, n132, n133, n136, n137, n138,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n153, n155, n156, n157, n158, n160, n163, n164, n165, n166,
         n167, n169, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n201, n203,
         n204, n205, n206, n207, n209, n211, n212, n213, n214, n215, n217,
         n219, n220, n221, n222, n223, n225, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n237, n239, n240, n241, n242, n243, n245,
         n247, n253, n254, n255, n256, n258, n259, n260, n263, n267, n268,
         n270, n271, n273, n276, n277, n278, n281, n282, n286, n290, n293,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438;

  AOI21X1 U17 ( .A0(n51), .A1(n68), .B0(n52), .Y(n50) );
  NOR2X2 U18 ( .A(n60), .B(n53), .Y(n51) );
  NOR2X2 U34 ( .A(B[36]), .B(A[36]), .Y(n60) );
  AOI21X1 U53 ( .A0(n86), .A1(n78), .B0(n79), .Y(n77) );
  AOI21X1 U77 ( .A0(n104), .A1(n96), .B0(n97), .Y(n95) );
  AOI21X1 U108 ( .A0(n131), .A1(n118), .B0(n119), .Y(n117) );
  AOI21X1 U116 ( .A0(n123), .A1(n143), .B0(n124), .Y(n122) );
  AOI21X1 U126 ( .A0(n143), .A1(n130), .B0(n131), .Y(n129) );
  AOI21X1 U138 ( .A0(n143), .A1(n270), .B0(n140), .Y(n138) );
  AOI21X1 U157 ( .A0(n430), .A1(n160), .B0(n153), .Y(n151) );
  AOI21X1 U315 ( .A0(n432), .A1(n427), .B0(n245), .Y(n243) );
  OAI21X2 U340 ( .A0(n173), .A1(n175), .B0(n174), .Y(n172) );
  NOR2X1 U341 ( .A(n91), .B(n98), .Y(n89) );
  AOI21X1 U342 ( .A0(n145), .A1(n164), .B0(n146), .Y(n144) );
  NOR2X1 U343 ( .A(n150), .B(n147), .Y(n145) );
  OAI21X1 U344 ( .A0(n151), .A1(n147), .B0(n148), .Y(n146) );
  OAI21X1 U345 ( .A0(n116), .A1(n144), .B0(n117), .Y(n115) );
  NAND2X1 U346 ( .A(n130), .B(n118), .Y(n116) );
  NOR2X1 U347 ( .A(n125), .B(n120), .Y(n118) );
  AOI21X1 U348 ( .A0(n89), .A1(n104), .B0(n90), .Y(n84) );
  NOR2X1 U349 ( .A(B[37]), .B(A[37]), .Y(n53) );
  OAI21X1 U350 ( .A0(n165), .A1(n167), .B0(n166), .Y(n164) );
  NOR2X1 U351 ( .A(B[25]), .B(A[25]), .Y(n147) );
  NOR2X1 U352 ( .A(B[29]), .B(A[29]), .Y(n120) );
  OAI21X1 U353 ( .A0(n142), .A1(n136), .B0(n137), .Y(n131) );
  NOR2X1 U354 ( .A(B[28]), .B(A[28]), .Y(n125) );
  NOR2X1 U355 ( .A(B[27]), .B(A[27]), .Y(n136) );
  INVX2 U356 ( .A(n115), .Y(n114) );
  NAND2X1 U357 ( .A(n67), .B(n51), .Y(n49) );
  NOR2X1 U358 ( .A(B[35]), .B(A[35]), .Y(n73) );
  OR2X1 U359 ( .A(n437), .B(A[39]), .Y(n426) );
  OAI21XL U360 ( .A0(n73), .A1(n81), .B0(n74), .Y(n68) );
  OAI21X1 U361 ( .A0(n84), .A1(n49), .B0(n50), .Y(n48) );
  NOR2X1 U362 ( .A(n49), .B(n83), .Y(n47) );
  INVX2 U363 ( .A(n84), .Y(n86) );
  OAI21X1 U364 ( .A0(n91), .A1(n99), .B0(n92), .Y(n90) );
  CLKINVX2 U365 ( .A(n83), .Y(n85) );
  INVXL U366 ( .A(n155), .Y(n153) );
  NOR2X1 U367 ( .A(B[19]), .B(A[19]), .Y(n178) );
  NOR2X1 U368 ( .A(B[31]), .B(A[31]), .Y(n109) );
  CLKINVXL U369 ( .A(n104), .Y(n102) );
  OAI21XL U370 ( .A0(n114), .A1(n65), .B0(n66), .Y(n64) );
  NAND2X1 U371 ( .A(n263), .B(n92), .Y(n7) );
  OAI21XL U372 ( .A0(n114), .A1(n56), .B0(n57), .Y(n55) );
  OAI21XL U373 ( .A0(n114), .A1(n76), .B0(n77), .Y(n75) );
  INVX1 U374 ( .A(n81), .Y(n79) );
  CLKINVX1 U375 ( .A(n158), .Y(n160) );
  OAI21XL U376 ( .A0(n53), .A1(n63), .B0(n54), .Y(n52) );
  INVX1 U377 ( .A(n44), .Y(n258) );
  NAND2BX1 U378 ( .AN(n73), .B(n74), .Y(n5) );
  NAND2XL U379 ( .A(n428), .B(n171), .Y(n19) );
  NOR2X1 U380 ( .A(B[26]), .B(A[26]), .Y(n141) );
  AOI21XL U381 ( .A0(n86), .A1(n67), .B0(n68), .Y(n66) );
  CLKINVXL U382 ( .A(n103), .Y(n101) );
  OAI21XL U383 ( .A0(n163), .A1(n150), .B0(n151), .Y(n149) );
  CLKINVXL U384 ( .A(n130), .Y(n132) );
  CLKINVXL U385 ( .A(n184), .Y(n183) );
  CLKINVXL U386 ( .A(n196), .Y(n195) );
  AOI21X1 U387 ( .A0(n58), .A1(n86), .B0(n59), .Y(n57) );
  NAND2X1 U388 ( .A(n58), .B(n85), .Y(n56) );
  OAI21X1 U389 ( .A0(n70), .A1(n60), .B0(n63), .Y(n59) );
  NAND2XL U390 ( .A(n260), .B(n63), .Y(n4) );
  CLKINVXL U391 ( .A(n99), .Y(n97) );
  NAND2XL U392 ( .A(n103), .B(n96), .Y(n94) );
  XOR2X1 U393 ( .A(n100), .B(n423), .Y(SUM[32]) );
  AND2X1 U394 ( .A(n96), .B(n99), .Y(n423) );
  NAND2XL U395 ( .A(n78), .B(n81), .Y(n6) );
  NAND2XL U396 ( .A(n267), .B(n121), .Y(n11) );
  NAND2XL U397 ( .A(n268), .B(n128), .Y(n12) );
  CLKINVXL U398 ( .A(n98), .Y(n96) );
  OAI21X2 U399 ( .A0(n109), .A1(n113), .B0(n110), .Y(n104) );
  NOR2BX1 U400 ( .AN(n67), .B(n60), .Y(n58) );
  NAND2XL U401 ( .A(n271), .B(n148), .Y(n15) );
  OAI21XL U402 ( .A0(n163), .A1(n157), .B0(n158), .Y(n156) );
  XOR2X1 U403 ( .A(n156), .B(n424), .Y(SUM[24]) );
  AND2X1 U404 ( .A(n430), .B(n155), .Y(n424) );
  CLKINVX2 U405 ( .A(n157), .Y(n273) );
  INVX1 U406 ( .A(n232), .Y(n231) );
  NAND2XL U407 ( .A(n276), .B(n174), .Y(n20) );
  NAND2XL U408 ( .A(n273), .B(n158), .Y(n17) );
  NAND2BXL U409 ( .AN(n109), .B(n110), .Y(n9) );
  CLKINVXL U410 ( .A(n173), .Y(n276) );
  XOR2X1 U411 ( .A(n180), .B(n425), .Y(SUM[19]) );
  AND2X1 U412 ( .A(n277), .B(n179), .Y(n425) );
  OAI21XL U413 ( .A0(n183), .A1(n181), .B0(n182), .Y(n180) );
  CLKINVXL U414 ( .A(n181), .Y(n278) );
  OAI21XL U415 ( .A0(n195), .A1(n193), .B0(n194), .Y(n192) );
  CLKINVXL U416 ( .A(n193), .Y(n281) );
  NAND2XL U417 ( .A(n282), .B(n198), .Y(n26) );
  CLKINVXL U418 ( .A(n197), .Y(n282) );
  NAND2XL U419 ( .A(n433), .B(n203), .Y(n27) );
  NAND2XL U420 ( .A(n435), .B(n211), .Y(n29) );
  NAND2XL U421 ( .A(n286), .B(n214), .Y(n30) );
  CLKINVXL U422 ( .A(n213), .Y(n286) );
  NAND2XL U423 ( .A(n434), .B(n219), .Y(n31) );
  NAND2XL U424 ( .A(n290), .B(n230), .Y(n34) );
  CLKINVXL U425 ( .A(n229), .Y(n290) );
  OR2XL U426 ( .A(B[24]), .B(A[24]), .Y(n430) );
  NAND2XL U427 ( .A(B[26]), .B(A[26]), .Y(n142) );
  NAND2XL U428 ( .A(B[30]), .B(A[30]), .Y(n113) );
  NOR2X1 U429 ( .A(B[33]), .B(A[33]), .Y(n91) );
  NAND2XL U430 ( .A(B[18]), .B(A[18]), .Y(n182) );
  NAND2XL U431 ( .A(B[15]), .B(A[15]), .Y(n194) );
  NAND2XL U432 ( .A(B[8]), .B(A[8]), .Y(n222) );
  OR2XL U433 ( .A(B[13]), .B(A[13]), .Y(n433) );
  NOR2X1 U434 ( .A(B[30]), .B(A[30]), .Y(n112) );
  NOR2XL U435 ( .A(B[34]), .B(A[34]), .Y(n80) );
  OR2XL U436 ( .A(B[7]), .B(A[7]), .Y(n431) );
  OR2XL U437 ( .A(B[21]), .B(A[21]), .Y(n428) );
  NAND2XL U438 ( .A(B[23]), .B(A[23]), .Y(n158) );
  NAND2XL U439 ( .A(B[21]), .B(A[21]), .Y(n171) );
  NAND2XL U440 ( .A(B[34]), .B(A[34]), .Y(n81) );
  NAND2XL U441 ( .A(B[7]), .B(A[7]), .Y(n227) );
  NAND2XL U442 ( .A(B[22]), .B(A[22]), .Y(n166) );
  NAND2X1 U443 ( .A(n426), .B(n42), .Y(n1) );
  NAND2XL U444 ( .A(n437), .B(A[38]), .Y(n45) );
  INVX2 U445 ( .A(n438), .Y(n437) );
  INVX2 U446 ( .A(B[38]), .Y(n438) );
  AOI21X1 U447 ( .A0(n115), .A1(n47), .B0(n48), .Y(n46) );
  INVX2 U448 ( .A(n68), .Y(n70) );
  OAI21XL U449 ( .A0(n114), .A1(n101), .B0(n102), .Y(n100) );
  OAI21XL U450 ( .A0(n114), .A1(n83), .B0(n84), .Y(n82) );
  NAND2X1 U451 ( .A(n89), .B(n103), .Y(n83) );
  INVX2 U452 ( .A(n144), .Y(n143) );
  INVX2 U453 ( .A(n164), .Y(n163) );
  OAI21X1 U454 ( .A0(n46), .A1(n44), .B0(n45), .Y(n43) );
  NOR2X1 U455 ( .A(n80), .B(n73), .Y(n67) );
  XNOR2X1 U456 ( .A(n55), .B(n3), .Y(SUM[37]) );
  NAND2X1 U457 ( .A(n259), .B(n54), .Y(n3) );
  XOR2X1 U458 ( .A(n46), .B(n2), .Y(SUM[38]) );
  NAND2X1 U459 ( .A(n258), .B(n45), .Y(n2) );
  XNOR2X1 U460 ( .A(n64), .B(n4), .Y(SUM[36]) );
  NOR2X1 U461 ( .A(n141), .B(n136), .Y(n130) );
  OAI21XL U462 ( .A0(n120), .A1(n128), .B0(n121), .Y(n119) );
  OAI21XL U463 ( .A0(n114), .A1(n94), .B0(n95), .Y(n93) );
  XNOR2X1 U464 ( .A(n93), .B(n7), .Y(SUM[33]) );
  OAI21XL U465 ( .A0(n114), .A1(n112), .B0(n113), .Y(n111) );
  XNOR2X1 U466 ( .A(n82), .B(n6), .Y(SUM[34]) );
  NAND2XL U467 ( .A(n85), .B(n78), .Y(n76) );
  AOI21X1 U468 ( .A0(n172), .A1(n428), .B0(n169), .Y(n167) );
  INVX2 U469 ( .A(n171), .Y(n169) );
  AOI21X1 U470 ( .A0(n176), .A1(n184), .B0(n177), .Y(n175) );
  OAI21X1 U471 ( .A0(n178), .A1(n182), .B0(n179), .Y(n177) );
  NOR2X1 U472 ( .A(n181), .B(n178), .Y(n176) );
  OAI21X1 U473 ( .A0(n213), .A1(n215), .B0(n214), .Y(n212) );
  OAI21X1 U474 ( .A0(n221), .A1(n223), .B0(n222), .Y(n220) );
  AOI21X1 U475 ( .A0(n204), .A1(n433), .B0(n201), .Y(n199) );
  INVX2 U476 ( .A(n203), .Y(n201) );
  AOI21X1 U477 ( .A0(n435), .A1(n212), .B0(n209), .Y(n207) );
  INVX2 U478 ( .A(n211), .Y(n209) );
  OAI21X1 U479 ( .A0(n199), .A1(n197), .B0(n198), .Y(n196) );
  AOI21X1 U480 ( .A0(n188), .A1(n196), .B0(n189), .Y(n187) );
  OAI21X1 U481 ( .A0(n190), .A1(n194), .B0(n191), .Y(n189) );
  NOR2X1 U482 ( .A(n193), .B(n190), .Y(n188) );
  OAI21X1 U483 ( .A0(n187), .A1(n185), .B0(n186), .Y(n184) );
  AOI21X1 U484 ( .A0(n220), .A1(n434), .B0(n217), .Y(n215) );
  INVX2 U485 ( .A(n219), .Y(n217) );
  OAI21X1 U486 ( .A0(n205), .A1(n207), .B0(n206), .Y(n204) );
  AOI21X1 U487 ( .A0(n429), .A1(n240), .B0(n237), .Y(n235) );
  INVX2 U488 ( .A(n239), .Y(n237) );
  OAI21X1 U489 ( .A0(n229), .A1(n231), .B0(n230), .Y(n228) );
  AOI21X1 U490 ( .A0(n228), .A1(n431), .B0(n225), .Y(n223) );
  INVX2 U491 ( .A(n227), .Y(n225) );
  OAI21X1 U492 ( .A0(n233), .A1(n235), .B0(n234), .Y(n232) );
  NOR2X1 U493 ( .A(n112), .B(n109), .Y(n103) );
  XOR2X1 U494 ( .A(n129), .B(n12), .Y(SUM[28]) );
  OAI21XL U495 ( .A0(n133), .A1(n125), .B0(n128), .Y(n124) );
  NOR2X1 U496 ( .A(n132), .B(n125), .Y(n123) );
  CLKINVXL U497 ( .A(n131), .Y(n133) );
  INVX2 U498 ( .A(n247), .Y(n245) );
  OAI21X1 U499 ( .A0(n241), .A1(n243), .B0(n242), .Y(n240) );
  INVX2 U500 ( .A(n142), .Y(n140) );
  NAND2X1 U501 ( .A(n273), .B(n430), .Y(n150) );
  INVX2 U502 ( .A(n80), .Y(n78) );
  CLKINVXL U503 ( .A(n60), .Y(n260) );
  CLKINVXL U504 ( .A(n53), .Y(n259) );
  OAI2BB1X1 U505 ( .A0N(n436), .A1N(n254), .B0(n253), .Y(n427) );
  XNOR2X1 U506 ( .A(n149), .B(n15), .Y(SUM[25]) );
  INVX2 U507 ( .A(n141), .Y(n270) );
  CLKINVXL U508 ( .A(n120), .Y(n267) );
  CLKINVXL U509 ( .A(n125), .Y(n268) );
  NAND2BX1 U510 ( .AN(n136), .B(n137), .Y(n13) );
  CLKINVXL U511 ( .A(n147), .Y(n271) );
  INVX2 U512 ( .A(n91), .Y(n263) );
  NAND2X1 U513 ( .A(n270), .B(n142), .Y(n14) );
  INVX2 U514 ( .A(n256), .Y(n254) );
  NAND2BX1 U515 ( .AN(n112), .B(n113), .Y(n10) );
  XOR2XL U516 ( .A(n20), .B(n175), .Y(SUM[20]) );
  NAND2BX1 U517 ( .AN(n165), .B(n166), .Y(n18) );
  XOR2X1 U518 ( .A(n183), .B(n22), .Y(SUM[18]) );
  NAND2X1 U519 ( .A(n278), .B(n182), .Y(n22) );
  NAND2BX1 U520 ( .AN(n185), .B(n186), .Y(n23) );
  INVX2 U521 ( .A(n178), .Y(n277) );
  XOR2X1 U522 ( .A(n25), .B(n195), .Y(SUM[15]) );
  NAND2X1 U523 ( .A(n281), .B(n194), .Y(n25) );
  NAND2BX1 U524 ( .AN(n190), .B(n191), .Y(n24) );
  XOR2XL U525 ( .A(n26), .B(n199), .Y(SUM[14]) );
  NAND2BX1 U526 ( .AN(n205), .B(n206), .Y(n28) );
  XNOR2XL U527 ( .A(n29), .B(n212), .Y(SUM[11]) );
  NAND2X1 U528 ( .A(n431), .B(n227), .Y(n33) );
  NAND2BX1 U529 ( .AN(n221), .B(n222), .Y(n32) );
  XOR2XL U530 ( .A(n34), .B(n231), .Y(SUM[6]) );
  NAND2XL U531 ( .A(n429), .B(n239), .Y(n36) );
  NAND2BX1 U532 ( .AN(n233), .B(n234), .Y(n35) );
  XOR2X1 U533 ( .A(n37), .B(n243), .Y(SUM[3]) );
  NAND2X1 U534 ( .A(n293), .B(n242), .Y(n37) );
  INVX2 U535 ( .A(n241), .Y(n293) );
  XNOR2X1 U536 ( .A(n38), .B(n427), .Y(SUM[2]) );
  NAND2X1 U537 ( .A(n432), .B(n247), .Y(n38) );
  NAND2X1 U538 ( .A(n436), .B(n253), .Y(n39) );
  XNOR2X1 U539 ( .A(n43), .B(n1), .Y(SUM[39]) );
  XNOR2X1 U540 ( .A(n111), .B(n9), .Y(SUM[31]) );
  XNOR2X1 U541 ( .A(n75), .B(n5), .Y(SUM[35]) );
  NOR2X1 U542 ( .A(B[20]), .B(A[20]), .Y(n173) );
  NOR2X1 U543 ( .A(B[18]), .B(A[18]), .Y(n181) );
  NAND2XL U544 ( .A(B[36]), .B(A[36]), .Y(n63) );
  NOR2X1 U545 ( .A(B[14]), .B(A[14]), .Y(n197) );
  NOR2X1 U546 ( .A(B[16]), .B(A[16]), .Y(n190) );
  NOR2X1 U547 ( .A(B[15]), .B(A[15]), .Y(n193) );
  NAND2XL U548 ( .A(B[35]), .B(A[35]), .Y(n74) );
  NAND2XL U549 ( .A(B[37]), .B(A[37]), .Y(n54) );
  NOR2X1 U550 ( .A(B[32]), .B(A[32]), .Y(n98) );
  XOR2X1 U551 ( .A(n114), .B(n10), .Y(SUM[30]) );
  NAND2XL U552 ( .A(B[20]), .B(A[20]), .Y(n174) );
  OR2XL U553 ( .A(B[4]), .B(A[4]), .Y(n429) );
  NOR2X1 U554 ( .A(B[17]), .B(A[17]), .Y(n185) );
  NAND2XL U555 ( .A(B[19]), .B(A[19]), .Y(n179) );
  NAND2XL U556 ( .A(B[27]), .B(A[27]), .Y(n137) );
  NAND2XL U557 ( .A(B[14]), .B(A[14]), .Y(n198) );
  NOR2X1 U558 ( .A(B[5]), .B(A[5]), .Y(n233) );
  NOR2X1 U559 ( .A(B[10]), .B(A[10]), .Y(n213) );
  NAND2XL U560 ( .A(B[28]), .B(A[28]), .Y(n128) );
  OR2XL U561 ( .A(B[2]), .B(A[2]), .Y(n432) );
  NOR2X1 U562 ( .A(B[12]), .B(A[12]), .Y(n205) );
  XOR2X1 U563 ( .A(n138), .B(n13), .Y(SUM[27]) );
  NAND2XL U564 ( .A(B[16]), .B(A[16]), .Y(n191) );
  NOR2X1 U565 ( .A(B[6]), .B(A[6]), .Y(n229) );
  OR2XL U566 ( .A(B[9]), .B(A[9]), .Y(n434) );
  NOR2X1 U567 ( .A(B[23]), .B(A[23]), .Y(n157) );
  NOR2X1 U568 ( .A(B[8]), .B(A[8]), .Y(n221) );
  NAND2XL U569 ( .A(B[29]), .B(A[29]), .Y(n121) );
  NAND2XL U570 ( .A(B[24]), .B(A[24]), .Y(n155) );
  OR2XL U571 ( .A(B[11]), .B(A[11]), .Y(n435) );
  NAND2XL U572 ( .A(B[13]), .B(A[13]), .Y(n203) );
  NOR2X1 U573 ( .A(n437), .B(A[38]), .Y(n44) );
  NAND2XL U574 ( .A(B[2]), .B(A[2]), .Y(n247) );
  NAND2XL U575 ( .A(B[17]), .B(A[17]), .Y(n186) );
  NAND2XL U576 ( .A(B[5]), .B(A[5]), .Y(n234) );
  NAND2XL U577 ( .A(B[9]), .B(A[9]), .Y(n219) );
  NAND2XL U578 ( .A(B[25]), .B(A[25]), .Y(n148) );
  OR2XL U579 ( .A(B[1]), .B(A[1]), .Y(n436) );
  NAND2XL U580 ( .A(B[33]), .B(A[33]), .Y(n92) );
  NAND2XL U581 ( .A(B[31]), .B(A[31]), .Y(n110) );
  NAND2XL U582 ( .A(B[12]), .B(A[12]), .Y(n206) );
  NAND2XL U583 ( .A(B[6]), .B(A[6]), .Y(n230) );
  NAND2XL U584 ( .A(B[10]), .B(A[10]), .Y(n214) );
  NAND2X1 U585 ( .A(B[32]), .B(A[32]), .Y(n99) );
  NAND2XL U586 ( .A(B[11]), .B(A[11]), .Y(n211) );
  NAND2XL U587 ( .A(B[1]), .B(A[1]), .Y(n253) );
  NOR2X1 U588 ( .A(B[3]), .B(A[3]), .Y(n241) );
  NOR2X1 U589 ( .A(B[22]), .B(A[22]), .Y(n165) );
  XNOR2X1 U590 ( .A(n143), .B(n14), .Y(SUM[26]) );
  NAND2XL U591 ( .A(B[3]), .B(A[3]), .Y(n242) );
  XOR2X1 U592 ( .A(n163), .B(n17), .Y(SUM[23]) );
  NAND2X1 U593 ( .A(B[0]), .B(A[0]), .Y(n256) );
  XOR2XL U594 ( .A(n18), .B(n167), .Y(SUM[22]) );
  XOR2X1 U595 ( .A(n187), .B(n23), .Y(SUM[17]) );
  XNOR2X1 U596 ( .A(n192), .B(n24), .Y(SUM[16]) );
  XOR2XL U597 ( .A(n28), .B(n207), .Y(SUM[12]) );
  XNOR2XL U598 ( .A(n31), .B(n220), .Y(SUM[9]) );
  XNOR2X1 U599 ( .A(n39), .B(n254), .Y(SUM[1]) );
  NAND2BX1 U600 ( .AN(n255), .B(n256), .Y(n40) );
  NOR2X1 U601 ( .A(B[0]), .B(A[0]), .Y(n255) );
  INVX2 U602 ( .A(n40), .Y(SUM[0]) );
  NAND2X1 U603 ( .A(n437), .B(A[39]), .Y(n42) );
  NAND2XL U604 ( .A(B[4]), .B(A[4]), .Y(n239) );
  XNOR2X1 U605 ( .A(n172), .B(n19), .Y(SUM[21]) );
  XNOR2XL U606 ( .A(n33), .B(n228), .Y(SUM[7]) );
  XNOR2XL U607 ( .A(n27), .B(n204), .Y(SUM[13]) );
  XOR2XL U608 ( .A(n35), .B(n235), .Y(SUM[5]) );
  NAND2XL U609 ( .A(n85), .B(n67), .Y(n65) );
  XOR2XL U610 ( .A(n30), .B(n215), .Y(SUM[10]) );
  XNOR2XL U611 ( .A(n36), .B(n240), .Y(SUM[4]) );
  XOR2X1 U612 ( .A(n122), .B(n11), .Y(SUM[29]) );
  XOR2XL U613 ( .A(n32), .B(n223), .Y(SUM[8]) );
endmodule


module MMSA_DW01_add_34 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n20, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n63,
         n64, n65, n66, n67, n68, n69, n70, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n128, n129, n130, n131, n132, n133, n136, n137,
         n138, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n153, n155, n156, n157, n158, n160, n163, n164, n165,
         n166, n167, n169, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n201,
         n203, n204, n205, n206, n207, n209, n211, n212, n213, n214, n215,
         n217, n219, n220, n221, n222, n223, n225, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n237, n239, n240, n241, n242, n243,
         n245, n247, n253, n254, n255, n256, n259, n260, n263, n267, n268,
         n270, n271, n273, n276, n277, n278, n281, n282, n286, n290, n293,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438;

  AOI21X1 U27 ( .A0(n58), .A1(n86), .B0(n59), .Y(n57) );
  AOI21X1 U39 ( .A0(n86), .A1(n67), .B0(n68), .Y(n66) );
  AOI21X1 U53 ( .A0(n86), .A1(n78), .B0(n79), .Y(n77) );
  AOI21X1 U77 ( .A0(n104), .A1(n96), .B0(n97), .Y(n95) );
  NOR2X2 U92 ( .A(n112), .B(n109), .Y(n103) );
  AOI21X1 U108 ( .A0(n131), .A1(n118), .B0(n119), .Y(n117) );
  AOI21X1 U126 ( .A0(n143), .A1(n130), .B0(n131), .Y(n129) );
  AOI21X1 U138 ( .A0(n143), .A1(n270), .B0(n140), .Y(n138) );
  AOI21X1 U157 ( .A0(n434), .A1(n160), .B0(n153), .Y(n151) );
  AOI21X1 U280 ( .A0(n228), .A1(n429), .B0(n225), .Y(n223) );
  AOI21X2 U340 ( .A0(n176), .A1(n184), .B0(n177), .Y(n175) );
  OAI21X4 U341 ( .A0(n187), .A1(n185), .B0(n186), .Y(n184) );
  INVX4 U342 ( .A(n115), .Y(n114) );
  AOI21X2 U343 ( .A0(n188), .A1(n196), .B0(n189), .Y(n187) );
  OAI21X2 U344 ( .A0(n116), .A1(n144), .B0(n117), .Y(n115) );
  OAI21X1 U345 ( .A0(n165), .A1(n167), .B0(n166), .Y(n164) );
  NOR2X1 U346 ( .A(n91), .B(n98), .Y(n89) );
  AOI21X1 U347 ( .A0(n145), .A1(n164), .B0(n146), .Y(n144) );
  AOI21X1 U348 ( .A0(n89), .A1(n104), .B0(n90), .Y(n84) );
  NOR2X1 U349 ( .A(B[14]), .B(A[14]), .Y(n197) );
  NOR2X1 U350 ( .A(B[19]), .B(A[19]), .Y(n178) );
  NOR2X1 U351 ( .A(B[18]), .B(A[18]), .Y(n181) );
  NOR2X1 U352 ( .A(B[29]), .B(A[29]), .Y(n120) );
  OAI21X1 U353 ( .A0(n199), .A1(n197), .B0(n198), .Y(n196) );
  NOR2X1 U354 ( .A(B[33]), .B(A[33]), .Y(n91) );
  AOI21X1 U355 ( .A0(n172), .A1(n431), .B0(n169), .Y(n167) );
  NOR2X1 U356 ( .A(B[27]), .B(A[27]), .Y(n136) );
  NOR2X1 U357 ( .A(B[30]), .B(A[30]), .Y(n112) );
  AOI21X1 U358 ( .A0(n115), .A1(n47), .B0(n48), .Y(n46) );
  INVXL U359 ( .A(n155), .Y(n153) );
  NAND2X1 U360 ( .A(n130), .B(n118), .Y(n116) );
  OAI21X1 U361 ( .A0(n84), .A1(n49), .B0(n50), .Y(n48) );
  INVX1 U362 ( .A(n67), .Y(n69) );
  AOI21X1 U363 ( .A0(n123), .A1(n143), .B0(n124), .Y(n122) );
  OAI21XL U364 ( .A0(n133), .A1(n125), .B0(n128), .Y(n124) );
  AOI21XL U365 ( .A0(n51), .A1(n68), .B0(n52), .Y(n50) );
  INVX2 U366 ( .A(n84), .Y(n86) );
  INVX1 U367 ( .A(n130), .Y(n132) );
  CLKINVXL U368 ( .A(n144), .Y(n143) );
  OAI21XL U369 ( .A0(n114), .A1(n56), .B0(n57), .Y(n55) );
  CLKINVX1 U370 ( .A(n158), .Y(n160) );
  NAND2BX1 U371 ( .AN(n73), .B(n74), .Y(n5) );
  CLKINVX2 U372 ( .A(n83), .Y(n85) );
  OAI21XL U373 ( .A0(n163), .A1(n150), .B0(n151), .Y(n149) );
  NAND2X1 U374 ( .A(n58), .B(n85), .Y(n56) );
  OAI21X1 U375 ( .A0(n142), .A1(n136), .B0(n137), .Y(n131) );
  CLKINVXL U376 ( .A(n99), .Y(n97) );
  OAI21X1 U377 ( .A0(n120), .A1(n128), .B0(n121), .Y(n119) );
  XOR2X1 U378 ( .A(n100), .B(n423), .Y(SUM[32]) );
  AND2X1 U379 ( .A(n96), .B(n99), .Y(n423) );
  NAND2XL U380 ( .A(n263), .B(n92), .Y(n7) );
  NAND2XL U381 ( .A(n267), .B(n121), .Y(n11) );
  NAND2XL U382 ( .A(n268), .B(n128), .Y(n12) );
  CLKINVXL U383 ( .A(n98), .Y(n96) );
  OAI21X2 U384 ( .A0(n109), .A1(n113), .B0(n110), .Y(n104) );
  OAI21XL U385 ( .A0(n163), .A1(n157), .B0(n158), .Y(n156) );
  XOR2X1 U386 ( .A(n156), .B(n424), .Y(SUM[24]) );
  AND2X1 U387 ( .A(n434), .B(n155), .Y(n424) );
  NAND2XL U388 ( .A(n271), .B(n148), .Y(n15) );
  CLKINVX2 U389 ( .A(n157), .Y(n273) );
  INVX1 U390 ( .A(n68), .Y(n70) );
  OAI21XL U391 ( .A0(n53), .A1(n63), .B0(n54), .Y(n52) );
  CLKINVXL U392 ( .A(n141), .Y(n270) );
  CLKINVXL U393 ( .A(n147), .Y(n271) );
  CLKINVXL U394 ( .A(n125), .Y(n268) );
  INVX1 U395 ( .A(n232), .Y(n231) );
  XOR2X1 U396 ( .A(n172), .B(n425), .Y(SUM[21]) );
  AND2X1 U397 ( .A(n431), .B(n171), .Y(n425) );
  CLKINVXL U398 ( .A(n60), .Y(n260) );
  CLKINVXL U399 ( .A(n53), .Y(n259) );
  NAND2XL U400 ( .A(n78), .B(n81), .Y(n6) );
  NAND2XL U401 ( .A(n276), .B(n174), .Y(n20) );
  NAND2XL U402 ( .A(n273), .B(n158), .Y(n17) );
  CLKINVXL U403 ( .A(n173), .Y(n276) );
  XOR2X1 U404 ( .A(n180), .B(n426), .Y(SUM[19]) );
  AND2X1 U405 ( .A(n277), .B(n179), .Y(n426) );
  OAI21XL U406 ( .A0(n195), .A1(n193), .B0(n194), .Y(n192) );
  CLKINVXL U407 ( .A(n193), .Y(n281) );
  NAND2XL U408 ( .A(n433), .B(n211), .Y(n29) );
  NAND2XL U409 ( .A(n286), .B(n214), .Y(n30) );
  CLKINVXL U410 ( .A(n213), .Y(n286) );
  NAND2XL U411 ( .A(n290), .B(n230), .Y(n34) );
  CLKINVXL U412 ( .A(n229), .Y(n290) );
  OR2XL U413 ( .A(B[24]), .B(A[24]), .Y(n434) );
  NAND2XL U414 ( .A(B[26]), .B(A[26]), .Y(n142) );
  NAND2XL U415 ( .A(B[30]), .B(A[30]), .Y(n113) );
  NAND2XL U416 ( .A(B[23]), .B(A[23]), .Y(n158) );
  NAND2XL U417 ( .A(B[18]), .B(A[18]), .Y(n182) );
  NOR2XL U418 ( .A(B[35]), .B(A[35]), .Y(n73) );
  NAND2XL U419 ( .A(B[15]), .B(A[15]), .Y(n194) );
  NAND2XL U420 ( .A(B[8]), .B(A[8]), .Y(n222) );
  OR2XL U421 ( .A(B[13]), .B(A[13]), .Y(n428) );
  NOR2XL U422 ( .A(B[34]), .B(A[34]), .Y(n80) );
  NAND2XL U423 ( .A(B[34]), .B(A[34]), .Y(n81) );
  OR2XL U424 ( .A(B[21]), .B(A[21]), .Y(n431) );
  NAND2XL U425 ( .A(B[13]), .B(A[13]), .Y(n203) );
  OR2XL U426 ( .A(B[7]), .B(A[7]), .Y(n429) );
  NAND2XL U427 ( .A(B[21]), .B(A[21]), .Y(n171) );
  NAND2XL U428 ( .A(B[11]), .B(A[11]), .Y(n211) );
  NAND2XL U429 ( .A(B[14]), .B(A[14]), .Y(n198) );
  NAND2XL U430 ( .A(B[7]), .B(A[7]), .Y(n227) );
  NAND2XL U431 ( .A(B[22]), .B(A[22]), .Y(n166) );
  NAND2XL U432 ( .A(B[36]), .B(A[36]), .Y(n63) );
  OR2XL U433 ( .A(B[4]), .B(A[4]), .Y(n430) );
  NAND2XL U434 ( .A(B[4]), .B(A[4]), .Y(n239) );
  NAND2BX1 U435 ( .AN(n41), .B(n42), .Y(n1) );
  INVX2 U436 ( .A(n438), .Y(n437) );
  INVX2 U437 ( .A(B[38]), .Y(n438) );
  NAND2X1 U438 ( .A(n67), .B(n51), .Y(n49) );
  OAI21X1 U439 ( .A0(n114), .A1(n65), .B0(n66), .Y(n64) );
  NAND2X1 U440 ( .A(n85), .B(n67), .Y(n65) );
  NAND2X1 U441 ( .A(n89), .B(n103), .Y(n83) );
  OAI21XL U442 ( .A0(n114), .A1(n101), .B0(n102), .Y(n100) );
  INVX2 U443 ( .A(n104), .Y(n102) );
  CLKINVXL U444 ( .A(n103), .Y(n101) );
  OAI21XL U445 ( .A0(n114), .A1(n83), .B0(n84), .Y(n82) );
  CLKINVXL U446 ( .A(n164), .Y(n163) );
  INVX2 U447 ( .A(n184), .Y(n183) );
  INVX2 U448 ( .A(n196), .Y(n195) );
  NOR2X1 U449 ( .A(n80), .B(n73), .Y(n67) );
  NOR2X1 U450 ( .A(n69), .B(n60), .Y(n58) );
  XNOR2X1 U451 ( .A(n55), .B(n3), .Y(SUM[37]) );
  NAND2X1 U452 ( .A(n259), .B(n54), .Y(n3) );
  NOR2X1 U453 ( .A(n60), .B(n53), .Y(n51) );
  OAI21X1 U454 ( .A0(n73), .A1(n81), .B0(n74), .Y(n68) );
  XNOR2X1 U455 ( .A(n64), .B(n4), .Y(SUM[36]) );
  NAND2X1 U456 ( .A(n260), .B(n63), .Y(n4) );
  OAI21X1 U457 ( .A0(n70), .A1(n60), .B0(n63), .Y(n59) );
  OAI21X1 U458 ( .A0(n91), .A1(n99), .B0(n92), .Y(n90) );
  OAI21X1 U459 ( .A0(n190), .A1(n194), .B0(n191), .Y(n189) );
  NOR2X1 U460 ( .A(n193), .B(n190), .Y(n188) );
  OAI21X1 U461 ( .A0(n178), .A1(n182), .B0(n179), .Y(n177) );
  NOR2X1 U462 ( .A(n181), .B(n178), .Y(n176) );
  OAI21X1 U463 ( .A0(n173), .A1(n175), .B0(n174), .Y(n172) );
  INVX2 U464 ( .A(n171), .Y(n169) );
  OAI21X1 U465 ( .A0(n151), .A1(n147), .B0(n148), .Y(n146) );
  NOR2X1 U466 ( .A(n150), .B(n147), .Y(n145) );
  XOR2X1 U467 ( .A(n129), .B(n12), .Y(SUM[28]) );
  NOR2X1 U468 ( .A(n141), .B(n136), .Y(n130) );
  OAI21XL U469 ( .A0(n114), .A1(n94), .B0(n95), .Y(n93) );
  NAND2XL U470 ( .A(n103), .B(n96), .Y(n94) );
  XNOR2X1 U471 ( .A(n93), .B(n7), .Y(SUM[33]) );
  NOR2X1 U472 ( .A(n125), .B(n120), .Y(n118) );
  INVX2 U473 ( .A(n142), .Y(n140) );
  OAI21XL U474 ( .A0(n114), .A1(n76), .B0(n77), .Y(n75) );
  NAND2XL U475 ( .A(n85), .B(n78), .Y(n76) );
  INVX2 U476 ( .A(n81), .Y(n79) );
  OAI21XL U477 ( .A0(n114), .A1(n112), .B0(n113), .Y(n111) );
  AOI21X1 U478 ( .A0(n204), .A1(n428), .B0(n201), .Y(n199) );
  INVX2 U479 ( .A(n203), .Y(n201) );
  OAI21X1 U480 ( .A0(n221), .A1(n223), .B0(n222), .Y(n220) );
  AOI21X1 U481 ( .A0(n220), .A1(n435), .B0(n217), .Y(n215) );
  OAI21X1 U482 ( .A0(n205), .A1(n207), .B0(n206), .Y(n204) );
  INVX2 U483 ( .A(n227), .Y(n225) );
  AOI21X1 U484 ( .A0(n433), .A1(n212), .B0(n209), .Y(n207) );
  INVX2 U485 ( .A(n211), .Y(n209) );
  OAI21X1 U486 ( .A0(n213), .A1(n215), .B0(n214), .Y(n212) );
  OAI21X1 U487 ( .A0(n229), .A1(n231), .B0(n230), .Y(n228) );
  OAI21X1 U488 ( .A0(n233), .A1(n235), .B0(n234), .Y(n232) );
  NOR2X1 U489 ( .A(n132), .B(n125), .Y(n123) );
  CLKINVXL U490 ( .A(n131), .Y(n133) );
  XOR2X1 U491 ( .A(n122), .B(n11), .Y(SUM[29]) );
  AOI21X1 U492 ( .A0(n430), .A1(n240), .B0(n237), .Y(n235) );
  INVX2 U493 ( .A(n239), .Y(n237) );
  AOI21X1 U494 ( .A0(n432), .A1(n427), .B0(n245), .Y(n243) );
  INVX2 U495 ( .A(n247), .Y(n245) );
  OAI21X1 U496 ( .A0(n241), .A1(n243), .B0(n242), .Y(n240) );
  OAI2BB1X1 U497 ( .A0N(n436), .A1N(n254), .B0(n253), .Y(n427) );
  INVX2 U498 ( .A(n80), .Y(n78) );
  NAND2BX1 U499 ( .AN(n44), .B(n45), .Y(n2) );
  NAND2X1 U500 ( .A(n273), .B(n434), .Y(n150) );
  XNOR2X1 U501 ( .A(n149), .B(n15), .Y(SUM[25]) );
  CLKINVXL U502 ( .A(n120), .Y(n267) );
  CLKINVXL U503 ( .A(n91), .Y(n263) );
  NAND2BX1 U504 ( .AN(n136), .B(n137), .Y(n13) );
  INVX2 U505 ( .A(n256), .Y(n254) );
  NAND2BX1 U506 ( .AN(n112), .B(n113), .Y(n10) );
  NAND2BX1 U507 ( .AN(n109), .B(n110), .Y(n9) );
  NAND2X1 U508 ( .A(n270), .B(n142), .Y(n14) );
  XOR2XL U509 ( .A(n20), .B(n175), .Y(SUM[20]) );
  NAND2BX1 U510 ( .AN(n165), .B(n166), .Y(n18) );
  OAI21XL U511 ( .A0(n183), .A1(n181), .B0(n182), .Y(n180) );
  XOR2X1 U512 ( .A(n183), .B(n22), .Y(SUM[18]) );
  NAND2X1 U513 ( .A(n278), .B(n182), .Y(n22) );
  CLKINVXL U514 ( .A(n181), .Y(n278) );
  CLKINVXL U515 ( .A(n178), .Y(n277) );
  NAND2BX1 U516 ( .AN(n185), .B(n186), .Y(n23) );
  XOR2X1 U517 ( .A(n25), .B(n195), .Y(SUM[15]) );
  NAND2X1 U518 ( .A(n281), .B(n194), .Y(n25) );
  NAND2BX1 U519 ( .AN(n190), .B(n191), .Y(n24) );
  CLKINVXL U520 ( .A(n197), .Y(n282) );
  XOR2XL U521 ( .A(n26), .B(n199), .Y(SUM[14]) );
  NAND2X1 U522 ( .A(n282), .B(n198), .Y(n26) );
  NAND2X1 U523 ( .A(n428), .B(n203), .Y(n27) );
  NAND2BX1 U524 ( .AN(n205), .B(n206), .Y(n28) );
  XNOR2XL U525 ( .A(n29), .B(n212), .Y(SUM[11]) );
  XOR2XL U526 ( .A(n30), .B(n215), .Y(SUM[10]) );
  NAND2XL U527 ( .A(n435), .B(n219), .Y(n31) );
  NAND2BX1 U528 ( .AN(n221), .B(n222), .Y(n32) );
  XNOR2XL U529 ( .A(n33), .B(n228), .Y(SUM[7]) );
  NAND2X1 U530 ( .A(n429), .B(n227), .Y(n33) );
  XOR2XL U531 ( .A(n34), .B(n231), .Y(SUM[6]) );
  NAND2BX1 U532 ( .AN(n233), .B(n234), .Y(n35) );
  NAND2X1 U533 ( .A(n430), .B(n239), .Y(n36) );
  INVX2 U534 ( .A(n241), .Y(n293) );
  XOR2X1 U535 ( .A(n37), .B(n243), .Y(SUM[3]) );
  NAND2X1 U536 ( .A(n293), .B(n242), .Y(n37) );
  XNOR2X1 U537 ( .A(n38), .B(n427), .Y(SUM[2]) );
  NAND2X1 U538 ( .A(n432), .B(n247), .Y(n38) );
  NAND2X1 U539 ( .A(n436), .B(n253), .Y(n39) );
  XNOR2X1 U540 ( .A(n43), .B(n1), .Y(SUM[39]) );
  NOR2X1 U541 ( .A(B[37]), .B(A[37]), .Y(n53) );
  NOR2X1 U542 ( .A(B[36]), .B(A[36]), .Y(n60) );
  NOR2X1 U543 ( .A(B[31]), .B(A[31]), .Y(n109) );
  NAND2XL U544 ( .A(B[35]), .B(A[35]), .Y(n74) );
  NAND2XL U545 ( .A(B[37]), .B(A[37]), .Y(n54) );
  NOR2X1 U546 ( .A(B[28]), .B(A[28]), .Y(n125) );
  XOR2X1 U547 ( .A(n138), .B(n13), .Y(SUM[27]) );
  XNOR2X1 U548 ( .A(n75), .B(n5), .Y(SUM[35]) );
  XNOR2X1 U549 ( .A(n111), .B(n9), .Y(SUM[31]) );
  XNOR2X1 U550 ( .A(n82), .B(n6), .Y(SUM[34]) );
  NOR2X1 U551 ( .A(B[16]), .B(A[16]), .Y(n190) );
  NOR2X1 U552 ( .A(B[20]), .B(A[20]), .Y(n173) );
  NOR2X1 U553 ( .A(B[26]), .B(A[26]), .Y(n141) );
  NOR2X1 U554 ( .A(B[5]), .B(A[5]), .Y(n233) );
  NOR2X1 U555 ( .A(B[32]), .B(A[32]), .Y(n98) );
  NOR2X1 U556 ( .A(B[15]), .B(A[15]), .Y(n193) );
  NOR2X1 U557 ( .A(B[6]), .B(A[6]), .Y(n229) );
  XOR2X1 U558 ( .A(n114), .B(n10), .Y(SUM[30]) );
  NOR2X1 U559 ( .A(B[12]), .B(A[12]), .Y(n205) );
  NOR2X1 U560 ( .A(B[17]), .B(A[17]), .Y(n185) );
  NOR2X1 U561 ( .A(B[25]), .B(A[25]), .Y(n147) );
  NOR2X1 U562 ( .A(B[10]), .B(A[10]), .Y(n213) );
  OR2XL U563 ( .A(B[2]), .B(A[2]), .Y(n432) );
  NAND2XL U564 ( .A(B[20]), .B(A[20]), .Y(n174) );
  OR2XL U565 ( .A(B[11]), .B(A[11]), .Y(n433) );
  NAND2XL U566 ( .A(B[27]), .B(A[27]), .Y(n137) );
  NAND2XL U567 ( .A(B[5]), .B(A[5]), .Y(n234) );
  NAND2XL U568 ( .A(B[19]), .B(A[19]), .Y(n179) );
  NOR2X1 U569 ( .A(n437), .B(A[38]), .Y(n44) );
  NOR2X1 U570 ( .A(B[3]), .B(A[3]), .Y(n241) );
  NAND2XL U571 ( .A(B[28]), .B(A[28]), .Y(n128) );
  NOR2X1 U572 ( .A(B[8]), .B(A[8]), .Y(n221) );
  NAND2XL U573 ( .A(B[16]), .B(A[16]), .Y(n191) );
  NAND2XL U574 ( .A(B[6]), .B(A[6]), .Y(n230) );
  OR2XL U575 ( .A(B[9]), .B(A[9]), .Y(n435) );
  NAND2XL U576 ( .A(B[33]), .B(A[33]), .Y(n92) );
  NAND2X1 U577 ( .A(B[32]), .B(A[32]), .Y(n99) );
  OR2XL U578 ( .A(B[1]), .B(A[1]), .Y(n436) );
  NAND2XL U579 ( .A(B[31]), .B(A[31]), .Y(n110) );
  NAND2XL U580 ( .A(B[2]), .B(A[2]), .Y(n247) );
  NAND2XL U581 ( .A(B[12]), .B(A[12]), .Y(n206) );
  NAND2XL U582 ( .A(B[29]), .B(A[29]), .Y(n121) );
  NOR2X1 U583 ( .A(B[23]), .B(A[23]), .Y(n157) );
  NAND2XL U584 ( .A(B[17]), .B(A[17]), .Y(n186) );
  NAND2XL U585 ( .A(B[24]), .B(A[24]), .Y(n155) );
  NAND2XL U586 ( .A(n437), .B(A[39]), .Y(n42) );
  NOR2X1 U587 ( .A(n437), .B(A[39]), .Y(n41) );
  NAND2XL U588 ( .A(n437), .B(A[38]), .Y(n45) );
  NAND2XL U589 ( .A(B[10]), .B(A[10]), .Y(n214) );
  NAND2XL U590 ( .A(B[25]), .B(A[25]), .Y(n148) );
  XNOR2X1 U591 ( .A(n143), .B(n14), .Y(SUM[26]) );
  NAND2XL U592 ( .A(B[1]), .B(A[1]), .Y(n253) );
  NAND2XL U593 ( .A(B[3]), .B(A[3]), .Y(n242) );
  NOR2X1 U594 ( .A(B[22]), .B(A[22]), .Y(n165) );
  XOR2X1 U595 ( .A(n163), .B(n17), .Y(SUM[23]) );
  NAND2X1 U596 ( .A(B[0]), .B(A[0]), .Y(n256) );
  XOR2XL U597 ( .A(n18), .B(n167), .Y(SUM[22]) );
  XNOR2X1 U598 ( .A(n192), .B(n24), .Y(SUM[16]) );
  XNOR2XL U599 ( .A(n27), .B(n204), .Y(SUM[13]) );
  XNOR2XL U600 ( .A(n31), .B(n220), .Y(SUM[9]) );
  XOR2XL U601 ( .A(n35), .B(n235), .Y(SUM[5]) );
  XNOR2XL U602 ( .A(n36), .B(n240), .Y(SUM[4]) );
  XNOR2X1 U603 ( .A(n39), .B(n254), .Y(SUM[1]) );
  NAND2BX1 U604 ( .AN(n255), .B(n256), .Y(n40) );
  NOR2X1 U605 ( .A(B[0]), .B(A[0]), .Y(n255) );
  INVX2 U606 ( .A(n40), .Y(SUM[0]) );
  INVX2 U607 ( .A(n219), .Y(n217) );
  NAND2XL U608 ( .A(B[9]), .B(A[9]), .Y(n219) );
  XOR2X1 U609 ( .A(n46), .B(n2), .Y(SUM[38]) );
  XOR2X1 U610 ( .A(n187), .B(n23), .Y(SUM[17]) );
  XOR2XL U611 ( .A(n32), .B(n223), .Y(SUM[8]) );
  XOR2XL U612 ( .A(n28), .B(n207), .Y(SUM[12]) );
  OAI21X1 U613 ( .A0(n46), .A1(n44), .B0(n45), .Y(n43) );
  NOR2X1 U614 ( .A(n49), .B(n83), .Y(n47) );
endmodule


module MMSA_DW01_add_33 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n7, n9, n10, n11, n12, n13, n14, n16, n17, n18,
         n20, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n63, n64,
         n65, n66, n67, n68, n69, n70, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n128, n129, n130, n131, n132, n133, n136, n137, n138,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n153, n155, n156, n157, n158, n160, n163, n164, n165, n166,
         n167, n169, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n201, n203,
         n204, n205, n206, n207, n209, n211, n212, n213, n214, n215, n217,
         n219, n220, n221, n222, n223, n225, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n237, n239, n240, n241, n242, n243, n245,
         n247, n253, n254, n255, n256, n258, n259, n260, n263, n267, n268,
         n270, n271, n273, n276, n277, n278, n281, n282, n286, n290, n293,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439;

  AOI21X1 U17 ( .A0(n51), .A1(n68), .B0(n52), .Y(n50) );
  AOI21X1 U27 ( .A0(n58), .A1(n86), .B0(n59), .Y(n57) );
  AOI21X1 U39 ( .A0(n86), .A1(n67), .B0(n68), .Y(n66) );
  AOI21X1 U53 ( .A0(n86), .A1(n78), .B0(n79), .Y(n77) );
  AOI21X1 U77 ( .A0(n104), .A1(n96), .B0(n97), .Y(n95) );
  AOI21X1 U108 ( .A0(n131), .A1(n118), .B0(n119), .Y(n117) );
  AOI21X1 U116 ( .A0(n123), .A1(n143), .B0(n124), .Y(n122) );
  AOI21X1 U126 ( .A0(n143), .A1(n130), .B0(n131), .Y(n129) );
  AOI21X1 U138 ( .A0(n143), .A1(n270), .B0(n140), .Y(n138) );
  AOI21X1 U157 ( .A0(n436), .A1(n160), .B0(n153), .Y(n151) );
  OAI21X1 U340 ( .A0(n165), .A1(n167), .B0(n166), .Y(n164) );
  AOI21X1 U341 ( .A0(n145), .A1(n164), .B0(n146), .Y(n144) );
  NOR2X1 U342 ( .A(B[14]), .B(A[14]), .Y(n197) );
  NOR2X1 U343 ( .A(B[19]), .B(A[19]), .Y(n178) );
  NOR2X1 U344 ( .A(B[18]), .B(A[18]), .Y(n181) );
  OAI21X1 U345 ( .A0(n116), .A1(n144), .B0(n117), .Y(n115) );
  NOR2X1 U346 ( .A(n80), .B(n73), .Y(n67) );
  NOR2X1 U347 ( .A(B[27]), .B(A[27]), .Y(n136) );
  INVX2 U348 ( .A(n115), .Y(n114) );
  OAI21XL U349 ( .A0(n114), .A1(n101), .B0(n102), .Y(n100) );
  INVXL U350 ( .A(n155), .Y(n153) );
  OAI21X1 U351 ( .A0(n73), .A1(n81), .B0(n74), .Y(n68) );
  CLKINVX2 U352 ( .A(n83), .Y(n85) );
  NOR2X1 U353 ( .A(B[33]), .B(A[33]), .Y(n91) );
  CLKINVXL U354 ( .A(n99), .Y(n97) );
  NOR2X1 U355 ( .A(n141), .B(n136), .Y(n130) );
  INVX1 U356 ( .A(n81), .Y(n79) );
  NAND2XL U357 ( .A(n436), .B(n155), .Y(n16) );
  INVX1 U358 ( .A(n44), .Y(n258) );
  NAND2XL U359 ( .A(n85), .B(n67), .Y(n65) );
  AOI21XL U360 ( .A0(n115), .A1(n47), .B0(n48), .Y(n46) );
  CLKINVXL U361 ( .A(n104), .Y(n102) );
  CLKINVXL U362 ( .A(n103), .Y(n101) );
  CLKINVXL U363 ( .A(n144), .Y(n143) );
  OAI21XL U364 ( .A0(n163), .A1(n150), .B0(n151), .Y(n149) );
  CLKINVXL U365 ( .A(n184), .Y(n183) );
  CLKINVXL U366 ( .A(n196), .Y(n195) );
  NAND2XL U367 ( .A(n103), .B(n96), .Y(n94) );
  CLKINVX1 U368 ( .A(n158), .Y(n160) );
  NAND2X1 U369 ( .A(n130), .B(n118), .Y(n116) );
  OAI21X1 U370 ( .A0(n120), .A1(n128), .B0(n121), .Y(n119) );
  OAI21X1 U371 ( .A0(n46), .A1(n44), .B0(n45), .Y(n43) );
  AOI21X1 U372 ( .A0(n89), .A1(n104), .B0(n90), .Y(n84) );
  OAI21XL U373 ( .A0(n91), .A1(n99), .B0(n92), .Y(n90) );
  XOR2X1 U374 ( .A(n100), .B(n423), .Y(SUM[32]) );
  AND2X1 U375 ( .A(n96), .B(n99), .Y(n423) );
  OAI21X1 U376 ( .A0(n142), .A1(n136), .B0(n137), .Y(n131) );
  NAND2XL U377 ( .A(n85), .B(n78), .Y(n76) );
  XOR2X1 U378 ( .A(n82), .B(n424), .Y(SUM[34]) );
  AND2X1 U379 ( .A(n78), .B(n81), .Y(n424) );
  OAI21X1 U380 ( .A0(n173), .A1(n175), .B0(n174), .Y(n172) );
  CLKINVXL U381 ( .A(n131), .Y(n133) );
  OAI21XL U382 ( .A0(n133), .A1(n125), .B0(n128), .Y(n124) );
  NAND2XL U383 ( .A(n267), .B(n121), .Y(n11) );
  NAND2XL U384 ( .A(n268), .B(n128), .Y(n12) );
  CLKINVXL U385 ( .A(n98), .Y(n96) );
  CLKINVX2 U386 ( .A(n157), .Y(n273) );
  OAI21XL U387 ( .A0(n163), .A1(n157), .B0(n158), .Y(n156) );
  XOR2X1 U388 ( .A(n149), .B(n425), .Y(SUM[25]) );
  AND2X1 U389 ( .A(n271), .B(n148), .Y(n425) );
  INVX1 U390 ( .A(n68), .Y(n70) );
  OAI21XL U391 ( .A0(n53), .A1(n63), .B0(n54), .Y(n52) );
  INVX1 U392 ( .A(n232), .Y(n231) );
  CLKINVXL U393 ( .A(n141), .Y(n270) );
  CLKINVXL U394 ( .A(n147), .Y(n271) );
  CLKINVXL U395 ( .A(n125), .Y(n268) );
  CLKINVXL U396 ( .A(n80), .Y(n78) );
  CLKINVXL U397 ( .A(n60), .Y(n260) );
  CLKINVXL U398 ( .A(n120), .Y(n267) );
  CLKINVXL U399 ( .A(n53), .Y(n259) );
  XOR2X1 U400 ( .A(n172), .B(n426), .Y(SUM[21]) );
  AND2X1 U401 ( .A(n430), .B(n171), .Y(n426) );
  NAND2XL U402 ( .A(n276), .B(n174), .Y(n20) );
  NAND2XL U403 ( .A(n273), .B(n158), .Y(n17) );
  CLKINVXL U404 ( .A(n173), .Y(n276) );
  XOR2X1 U405 ( .A(n180), .B(n427), .Y(SUM[19]) );
  AND2X1 U406 ( .A(n277), .B(n179), .Y(n427) );
  OAI21XL U407 ( .A0(n195), .A1(n193), .B0(n194), .Y(n192) );
  CLKINVXL U408 ( .A(n193), .Y(n281) );
  NAND2XL U409 ( .A(n282), .B(n198), .Y(n26) );
  NAND2XL U410 ( .A(n434), .B(n203), .Y(n27) );
  NAND2XL U411 ( .A(n435), .B(n211), .Y(n29) );
  NAND2XL U412 ( .A(n286), .B(n214), .Y(n30) );
  CLKINVXL U413 ( .A(n213), .Y(n286) );
  NAND2XL U414 ( .A(n432), .B(n219), .Y(n31) );
  NAND2XL U415 ( .A(n290), .B(n230), .Y(n34) );
  CLKINVXL U416 ( .A(n229), .Y(n290) );
  OR2XL U417 ( .A(B[24]), .B(A[24]), .Y(n436) );
  NAND2XL U418 ( .A(B[24]), .B(A[24]), .Y(n155) );
  NAND2XL U419 ( .A(B[26]), .B(A[26]), .Y(n142) );
  NAND2XL U420 ( .A(B[18]), .B(A[18]), .Y(n182) );
  NAND2XL U421 ( .A(B[15]), .B(A[15]), .Y(n194) );
  NAND2XL U422 ( .A(B[8]), .B(A[8]), .Y(n222) );
  NAND2XL U423 ( .A(B[30]), .B(A[30]), .Y(n113) );
  OR2XL U424 ( .A(B[21]), .B(A[21]), .Y(n430) );
  OR2XL U425 ( .A(B[7]), .B(A[7]), .Y(n431) );
  NAND2XL U426 ( .A(B[21]), .B(A[21]), .Y(n171) );
  NAND2XL U427 ( .A(B[7]), .B(A[7]), .Y(n227) );
  NOR2X1 U428 ( .A(B[30]), .B(A[30]), .Y(n112) );
  NAND2XL U429 ( .A(B[34]), .B(A[34]), .Y(n81) );
  NAND2XL U430 ( .A(B[22]), .B(A[22]), .Y(n166) );
  NAND2XL U431 ( .A(B[36]), .B(A[36]), .Y(n63) );
  OR2XL U432 ( .A(B[4]), .B(A[4]), .Y(n429) );
  NAND2XL U433 ( .A(B[4]), .B(A[4]), .Y(n239) );
  NAND2BX1 U434 ( .AN(n41), .B(n42), .Y(n1) );
  NAND2XL U435 ( .A(n438), .B(A[38]), .Y(n45) );
  INVX2 U436 ( .A(n439), .Y(n438) );
  INVX2 U437 ( .A(B[38]), .Y(n439) );
  OAI21X1 U438 ( .A0(n84), .A1(n49), .B0(n50), .Y(n48) );
  NAND2X1 U439 ( .A(n67), .B(n51), .Y(n49) );
  INVX2 U440 ( .A(n67), .Y(n69) );
  OAI21XL U441 ( .A0(n114), .A1(n65), .B0(n66), .Y(n64) );
  OAI21XL U442 ( .A0(n114), .A1(n83), .B0(n84), .Y(n82) );
  NAND2X1 U443 ( .A(n89), .B(n103), .Y(n83) );
  INVX2 U444 ( .A(n84), .Y(n86) );
  INVX2 U445 ( .A(n130), .Y(n132) );
  CLKINVXL U446 ( .A(n164), .Y(n163) );
  NOR2X1 U447 ( .A(n60), .B(n53), .Y(n51) );
  OAI21XL U448 ( .A0(n114), .A1(n56), .B0(n57), .Y(n55) );
  NAND2X1 U449 ( .A(n58), .B(n85), .Y(n56) );
  NOR2X1 U450 ( .A(n69), .B(n60), .Y(n58) );
  XNOR2X1 U451 ( .A(n55), .B(n3), .Y(SUM[37]) );
  NAND2X1 U452 ( .A(n259), .B(n54), .Y(n3) );
  OAI21X1 U453 ( .A0(n70), .A1(n60), .B0(n63), .Y(n59) );
  NAND2X1 U454 ( .A(n258), .B(n45), .Y(n2) );
  NOR2X1 U455 ( .A(n132), .B(n125), .Y(n123) );
  AOI21X1 U456 ( .A0(n176), .A1(n184), .B0(n177), .Y(n175) );
  OAI21X1 U457 ( .A0(n178), .A1(n182), .B0(n179), .Y(n177) );
  NOR2X1 U458 ( .A(n181), .B(n178), .Y(n176) );
  AOI21X1 U459 ( .A0(n172), .A1(n430), .B0(n169), .Y(n167) );
  INVX2 U460 ( .A(n171), .Y(n169) );
  OAI21X1 U461 ( .A0(n151), .A1(n147), .B0(n148), .Y(n146) );
  NOR2X1 U462 ( .A(n150), .B(n147), .Y(n145) );
  XOR2X1 U463 ( .A(n122), .B(n11), .Y(SUM[29]) );
  OAI21XL U464 ( .A0(n114), .A1(n94), .B0(n95), .Y(n93) );
  XNOR2X1 U465 ( .A(n93), .B(n7), .Y(SUM[33]) );
  NAND2X1 U466 ( .A(n263), .B(n92), .Y(n7) );
  XNOR2X1 U467 ( .A(n64), .B(n4), .Y(SUM[36]) );
  NAND2X1 U468 ( .A(n260), .B(n63), .Y(n4) );
  XOR2X1 U469 ( .A(n129), .B(n12), .Y(SUM[28]) );
  OAI21X1 U470 ( .A0(n199), .A1(n197), .B0(n198), .Y(n196) );
  AOI21X1 U471 ( .A0(n188), .A1(n196), .B0(n189), .Y(n187) );
  OAI21X1 U472 ( .A0(n190), .A1(n194), .B0(n191), .Y(n189) );
  NOR2X1 U473 ( .A(n193), .B(n190), .Y(n188) );
  OAI21X1 U474 ( .A0(n187), .A1(n185), .B0(n186), .Y(n184) );
  OAI21XL U475 ( .A0(n114), .A1(n112), .B0(n113), .Y(n111) );
  OAI21XL U476 ( .A0(n114), .A1(n76), .B0(n77), .Y(n75) );
  AOI21X1 U477 ( .A0(n220), .A1(n432), .B0(n217), .Y(n215) );
  INVX2 U478 ( .A(n219), .Y(n217) );
  OAI21X1 U479 ( .A0(n205), .A1(n207), .B0(n206), .Y(n204) );
  AOI21X1 U480 ( .A0(n429), .A1(n240), .B0(n237), .Y(n235) );
  INVX2 U481 ( .A(n239), .Y(n237) );
  OAI21X1 U482 ( .A0(n213), .A1(n215), .B0(n214), .Y(n212) );
  OAI21X1 U483 ( .A0(n229), .A1(n231), .B0(n230), .Y(n228) );
  AOI21X1 U484 ( .A0(n435), .A1(n212), .B0(n209), .Y(n207) );
  INVX2 U485 ( .A(n211), .Y(n209) );
  OAI21X1 U486 ( .A0(n221), .A1(n223), .B0(n222), .Y(n220) );
  AOI21X1 U487 ( .A0(n204), .A1(n434), .B0(n201), .Y(n199) );
  INVX2 U488 ( .A(n203), .Y(n201) );
  AOI21X1 U489 ( .A0(n228), .A1(n431), .B0(n225), .Y(n223) );
  INVX2 U490 ( .A(n227), .Y(n225) );
  OAI21X1 U491 ( .A0(n233), .A1(n235), .B0(n234), .Y(n232) );
  INVX2 U492 ( .A(n142), .Y(n140) );
  NOR2X1 U493 ( .A(n125), .B(n120), .Y(n118) );
  NOR2X1 U494 ( .A(n91), .B(n98), .Y(n89) );
  OAI21X1 U495 ( .A0(n109), .A1(n113), .B0(n110), .Y(n104) );
  AOI21X1 U496 ( .A0(n433), .A1(n428), .B0(n245), .Y(n243) );
  INVX2 U497 ( .A(n247), .Y(n245) );
  OAI21X1 U498 ( .A0(n241), .A1(n243), .B0(n242), .Y(n240) );
  NOR2X1 U499 ( .A(n112), .B(n109), .Y(n103) );
  NAND2X1 U500 ( .A(n273), .B(n436), .Y(n150) );
  OAI2BB1X1 U501 ( .A0N(n437), .A1N(n254), .B0(n253), .Y(n428) );
  NAND2BX1 U502 ( .AN(n73), .B(n74), .Y(n5) );
  XNOR2X1 U503 ( .A(n156), .B(n16), .Y(SUM[24]) );
  NAND2BX1 U504 ( .AN(n136), .B(n137), .Y(n13) );
  INVX2 U505 ( .A(n256), .Y(n254) );
  INVX2 U506 ( .A(n91), .Y(n263) );
  NAND2X1 U507 ( .A(n270), .B(n142), .Y(n14) );
  NAND2BX1 U508 ( .AN(n112), .B(n113), .Y(n10) );
  NAND2BX1 U509 ( .AN(n109), .B(n110), .Y(n9) );
  XOR2XL U510 ( .A(n20), .B(n175), .Y(SUM[20]) );
  OAI21XL U511 ( .A0(n183), .A1(n181), .B0(n182), .Y(n180) );
  NAND2BX1 U512 ( .AN(n165), .B(n166), .Y(n18) );
  XOR2X1 U513 ( .A(n183), .B(n22), .Y(SUM[18]) );
  NAND2X1 U514 ( .A(n278), .B(n182), .Y(n22) );
  CLKINVXL U515 ( .A(n181), .Y(n278) );
  CLKINVXL U516 ( .A(n178), .Y(n277) );
  NAND2BX1 U517 ( .AN(n185), .B(n186), .Y(n23) );
  XOR2X1 U518 ( .A(n25), .B(n195), .Y(SUM[15]) );
  NAND2X1 U519 ( .A(n281), .B(n194), .Y(n25) );
  CLKINVXL U520 ( .A(n197), .Y(n282) );
  NAND2BX1 U521 ( .AN(n190), .B(n191), .Y(n24) );
  NAND2BX1 U522 ( .AN(n205), .B(n206), .Y(n28) );
  XNOR2XL U523 ( .A(n29), .B(n212), .Y(SUM[11]) );
  XOR2XL U524 ( .A(n30), .B(n215), .Y(SUM[10]) );
  NAND2BX1 U525 ( .AN(n221), .B(n222), .Y(n32) );
  XNOR2XL U526 ( .A(n33), .B(n228), .Y(SUM[7]) );
  NAND2X1 U527 ( .A(n431), .B(n227), .Y(n33) );
  XOR2XL U528 ( .A(n34), .B(n231), .Y(SUM[6]) );
  NAND2BX1 U529 ( .AN(n233), .B(n234), .Y(n35) );
  NAND2X1 U530 ( .A(n429), .B(n239), .Y(n36) );
  INVX2 U531 ( .A(n241), .Y(n293) );
  XOR2XL U532 ( .A(n37), .B(n243), .Y(SUM[3]) );
  NAND2X1 U533 ( .A(n293), .B(n242), .Y(n37) );
  XNOR2X1 U534 ( .A(n38), .B(n428), .Y(SUM[2]) );
  NAND2X1 U535 ( .A(n433), .B(n247), .Y(n38) );
  NAND2X1 U536 ( .A(n437), .B(n253), .Y(n39) );
  XNOR2X1 U537 ( .A(n43), .B(n1), .Y(SUM[39]) );
  NOR2X1 U538 ( .A(B[37]), .B(A[37]), .Y(n53) );
  NOR2X1 U539 ( .A(B[36]), .B(A[36]), .Y(n60) );
  NOR2X1 U540 ( .A(B[34]), .B(A[34]), .Y(n80) );
  NOR2X1 U541 ( .A(B[35]), .B(A[35]), .Y(n73) );
  NAND2XL U542 ( .A(B[35]), .B(A[35]), .Y(n74) );
  NAND2XL U543 ( .A(B[37]), .B(A[37]), .Y(n54) );
  NOR2X1 U544 ( .A(B[20]), .B(A[20]), .Y(n173) );
  XNOR2X1 U545 ( .A(n111), .B(n9), .Y(SUM[31]) );
  XNOR2X1 U546 ( .A(n75), .B(n5), .Y(SUM[35]) );
  NOR2X1 U547 ( .A(B[16]), .B(A[16]), .Y(n190) );
  XOR2X1 U548 ( .A(n138), .B(n13), .Y(SUM[27]) );
  NOR2X1 U549 ( .A(B[28]), .B(A[28]), .Y(n125) );
  NOR2X1 U550 ( .A(B[26]), .B(A[26]), .Y(n141) );
  NOR2X1 U551 ( .A(B[12]), .B(A[12]), .Y(n205) );
  NOR2X1 U552 ( .A(B[5]), .B(A[5]), .Y(n233) );
  NOR2X1 U553 ( .A(B[32]), .B(A[32]), .Y(n98) );
  NOR2X1 U554 ( .A(B[15]), .B(A[15]), .Y(n193) );
  NOR2X1 U555 ( .A(B[29]), .B(A[29]), .Y(n120) );
  XOR2X1 U556 ( .A(n114), .B(n10), .Y(SUM[30]) );
  NOR2X1 U557 ( .A(B[6]), .B(A[6]), .Y(n229) );
  NOR2X1 U558 ( .A(B[25]), .B(A[25]), .Y(n147) );
  NAND2X1 U559 ( .A(B[23]), .B(A[23]), .Y(n158) );
  OR2XL U560 ( .A(B[9]), .B(A[9]), .Y(n432) );
  NOR2X1 U561 ( .A(B[17]), .B(A[17]), .Y(n185) );
  NAND2XL U562 ( .A(B[28]), .B(A[28]), .Y(n128) );
  NOR2X1 U563 ( .A(B[31]), .B(A[31]), .Y(n109) );
  OR2XL U564 ( .A(B[2]), .B(A[2]), .Y(n433) );
  NOR2X1 U565 ( .A(B[10]), .B(A[10]), .Y(n213) );
  NAND2XL U566 ( .A(B[20]), .B(A[20]), .Y(n174) );
  OR2XL U567 ( .A(B[13]), .B(A[13]), .Y(n434) );
  OR2XL U568 ( .A(B[11]), .B(A[11]), .Y(n435) );
  NAND2XL U569 ( .A(B[19]), .B(A[19]), .Y(n179) );
  NAND2XL U570 ( .A(B[14]), .B(A[14]), .Y(n198) );
  NAND2XL U571 ( .A(B[27]), .B(A[27]), .Y(n137) );
  NAND2XL U572 ( .A(B[5]), .B(A[5]), .Y(n234) );
  NAND2XL U573 ( .A(B[9]), .B(A[9]), .Y(n219) );
  NOR2X1 U574 ( .A(n438), .B(A[38]), .Y(n44) );
  NOR2X1 U575 ( .A(B[8]), .B(A[8]), .Y(n221) );
  NAND2XL U576 ( .A(B[29]), .B(A[29]), .Y(n121) );
  NAND2XL U577 ( .A(B[11]), .B(A[11]), .Y(n211) );
  NOR2X1 U578 ( .A(B[3]), .B(A[3]), .Y(n241) );
  NAND2XL U579 ( .A(B[12]), .B(A[12]), .Y(n206) );
  NAND2XL U580 ( .A(B[33]), .B(A[33]), .Y(n92) );
  NAND2XL U581 ( .A(B[31]), .B(A[31]), .Y(n110) );
  NOR2X1 U582 ( .A(B[23]), .B(A[23]), .Y(n157) );
  NAND2XL U583 ( .A(B[16]), .B(A[16]), .Y(n191) );
  NAND2X1 U584 ( .A(B[32]), .B(A[32]), .Y(n99) );
  NAND2XL U585 ( .A(B[2]), .B(A[2]), .Y(n247) );
  NAND2XL U586 ( .A(B[6]), .B(A[6]), .Y(n230) );
  OR2XL U587 ( .A(B[1]), .B(A[1]), .Y(n437) );
  NAND2XL U588 ( .A(B[10]), .B(A[10]), .Y(n214) );
  NAND2XL U589 ( .A(B[13]), .B(A[13]), .Y(n203) );
  NAND2XL U590 ( .A(B[17]), .B(A[17]), .Y(n186) );
  NAND2X1 U591 ( .A(n438), .B(A[39]), .Y(n42) );
  NOR2X1 U592 ( .A(n438), .B(A[39]), .Y(n41) );
  NAND2XL U593 ( .A(B[25]), .B(A[25]), .Y(n148) );
  XNOR2X1 U594 ( .A(n143), .B(n14), .Y(SUM[26]) );
  NAND2XL U595 ( .A(B[1]), .B(A[1]), .Y(n253) );
  NAND2XL U596 ( .A(B[3]), .B(A[3]), .Y(n242) );
  NOR2X1 U597 ( .A(B[22]), .B(A[22]), .Y(n165) );
  XOR2X1 U598 ( .A(n163), .B(n17), .Y(SUM[23]) );
  NAND2X1 U599 ( .A(B[0]), .B(A[0]), .Y(n256) );
  XOR2XL U600 ( .A(n18), .B(n167), .Y(SUM[22]) );
  XOR2X1 U601 ( .A(n187), .B(n23), .Y(SUM[17]) );
  XNOR2X1 U602 ( .A(n192), .B(n24), .Y(SUM[16]) );
  XNOR2XL U603 ( .A(n27), .B(n204), .Y(SUM[13]) );
  XOR2XL U604 ( .A(n28), .B(n207), .Y(SUM[12]) );
  XNOR2XL U605 ( .A(n31), .B(n220), .Y(SUM[9]) );
  XOR2XL U606 ( .A(n35), .B(n235), .Y(SUM[5]) );
  XNOR2XL U607 ( .A(n36), .B(n240), .Y(SUM[4]) );
  XNOR2X1 U608 ( .A(n39), .B(n254), .Y(SUM[1]) );
  NAND2BX1 U609 ( .AN(n255), .B(n256), .Y(n40) );
  NOR2X1 U610 ( .A(B[0]), .B(A[0]), .Y(n255) );
  INVX2 U611 ( .A(n40), .Y(SUM[0]) );
  XOR2X1 U612 ( .A(n46), .B(n2), .Y(SUM[38]) );
  XOR2XL U613 ( .A(n26), .B(n199), .Y(SUM[14]) );
  XOR2XL U614 ( .A(n32), .B(n223), .Y(SUM[8]) );
  NOR2X1 U615 ( .A(n49), .B(n83), .Y(n47) );
endmodule


module MMSA_DW01_add_32 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n63, n64,
         n65, n66, n67, n68, n69, n70, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n128, n129, n130, n131, n132, n133, n136, n137, n138,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n153, n155, n156, n157, n158, n160, n163, n164, n165, n166,
         n167, n169, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n201, n203,
         n204, n205, n206, n207, n209, n211, n212, n213, n214, n215, n217,
         n219, n220, n221, n222, n223, n225, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n237, n239, n240, n241, n242, n243, n245,
         n247, n253, n254, n255, n256, n258, n259, n260, n263, n267, n268,
         n270, n271, n273, n276, n277, n278, n281, n282, n286, n290, n293,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438;

  AOI21X1 U13 ( .A0(n115), .A1(n47), .B0(n48), .Y(n46) );
  AOI21X1 U17 ( .A0(n51), .A1(n68), .B0(n52), .Y(n50) );
  AOI21X1 U27 ( .A0(n58), .A1(n86), .B0(n59), .Y(n57) );
  AOI21X1 U39 ( .A0(n86), .A1(n67), .B0(n68), .Y(n66) );
  AOI21X1 U53 ( .A0(n86), .A1(n78), .B0(n79), .Y(n77) );
  AOI21X1 U77 ( .A0(n104), .A1(n96), .B0(n97), .Y(n95) );
  AOI21X1 U108 ( .A0(n131), .A1(n118), .B0(n119), .Y(n117) );
  NOR2X2 U113 ( .A(B[29]), .B(A[29]), .Y(n120) );
  NOR2X2 U123 ( .A(B[28]), .B(A[28]), .Y(n125) );
  AOI21X1 U126 ( .A0(n143), .A1(n130), .B0(n131), .Y(n129) );
  AOI21X1 U138 ( .A0(n143), .A1(n270), .B0(n140), .Y(n138) );
  AOI21X1 U157 ( .A0(n429), .A1(n160), .B0(n153), .Y(n151) );
  AOI21X1 U196 ( .A0(n176), .A1(n184), .B0(n177), .Y(n175) );
  AOI21X1 U238 ( .A0(n204), .A1(n431), .B0(n201), .Y(n199) );
  AOI21X1 U266 ( .A0(n220), .A1(n428), .B0(n217), .Y(n215) );
  AOI21X1 U280 ( .A0(n228), .A1(n433), .B0(n225), .Y(n223) );
  AOI21X1 U301 ( .A0(n430), .A1(n240), .B0(n237), .Y(n235) );
  AOI21X1 U315 ( .A0(n434), .A1(n427), .B0(n245), .Y(n243) );
  NOR2XL U340 ( .A(B[35]), .B(A[35]), .Y(n73) );
  NOR2X1 U341 ( .A(B[19]), .B(A[19]), .Y(n178) );
  NOR2X1 U342 ( .A(B[18]), .B(A[18]), .Y(n181) );
  NOR2X1 U343 ( .A(B[16]), .B(A[16]), .Y(n190) );
  OAI21X1 U344 ( .A0(n116), .A1(n144), .B0(n117), .Y(n115) );
  NOR2X1 U345 ( .A(n80), .B(n73), .Y(n67) );
  NOR2X1 U346 ( .A(n112), .B(n109), .Y(n103) );
  NOR2X1 U347 ( .A(B[30]), .B(A[30]), .Y(n112) );
  INVX2 U348 ( .A(n115), .Y(n114) );
  OAI21X1 U349 ( .A0(n114), .A1(n101), .B0(n102), .Y(n100) );
  AOI21X2 U350 ( .A0(n145), .A1(n164), .B0(n146), .Y(n144) );
  OAI21X2 U351 ( .A0(n165), .A1(n167), .B0(n166), .Y(n164) );
  INVX2 U352 ( .A(n84), .Y(n86) );
  INVX1 U353 ( .A(n155), .Y(n153) );
  NOR2X1 U354 ( .A(B[27]), .B(A[27]), .Y(n136) );
  INVXL U355 ( .A(n103), .Y(n101) );
  NAND2X1 U356 ( .A(n89), .B(n103), .Y(n83) );
  NAND2X1 U357 ( .A(n58), .B(n85), .Y(n56) );
  OAI21X1 U358 ( .A0(n151), .A1(n147), .B0(n148), .Y(n146) );
  NAND2XL U359 ( .A(n78), .B(n81), .Y(n6) );
  CLKINVXL U360 ( .A(n81), .Y(n79) );
  CLKINVX1 U361 ( .A(n158), .Y(n160) );
  OAI21X1 U362 ( .A0(n70), .A1(n60), .B0(n63), .Y(n59) );
  INVX1 U363 ( .A(n44), .Y(n258) );
  OR2XL U364 ( .A(B[11]), .B(A[11]), .Y(n435) );
  CLKINVXL U365 ( .A(n104), .Y(n102) );
  OAI21XL U366 ( .A0(n114), .A1(n65), .B0(n66), .Y(n64) );
  OAI21XL U367 ( .A0(n163), .A1(n150), .B0(n151), .Y(n149) );
  CLKINVXL U368 ( .A(n164), .Y(n163) );
  CLKINVXL U369 ( .A(n184), .Y(n183) );
  CLKINVXL U370 ( .A(n196), .Y(n195) );
  CLKINVXL U371 ( .A(n99), .Y(n97) );
  NAND2XL U372 ( .A(n263), .B(n92), .Y(n7) );
  NAND2XL U373 ( .A(n96), .B(n99), .Y(n8) );
  AOI21X1 U374 ( .A0(n123), .A1(n143), .B0(n124), .Y(n122) );
  NAND2XL U375 ( .A(n267), .B(n121), .Y(n11) );
  NAND2XL U376 ( .A(n85), .B(n78), .Y(n76) );
  NAND2XL U377 ( .A(n268), .B(n128), .Y(n12) );
  CLKINVXL U378 ( .A(n142), .Y(n140) );
  CLKINVX1 U379 ( .A(n219), .Y(n217) );
  NOR2X2 U380 ( .A(n141), .B(n136), .Y(n130) );
  CLKINVX2 U381 ( .A(n157), .Y(n273) );
  NAND2XL U382 ( .A(n271), .B(n148), .Y(n15) );
  INVX1 U383 ( .A(n68), .Y(n70) );
  OAI21XL U384 ( .A0(n53), .A1(n63), .B0(n54), .Y(n52) );
  XOR2X1 U385 ( .A(n156), .B(n423), .Y(SUM[24]) );
  AND2X1 U386 ( .A(n429), .B(n155), .Y(n423) );
  OAI21XL U387 ( .A0(n163), .A1(n157), .B0(n158), .Y(n156) );
  INVX1 U388 ( .A(n232), .Y(n231) );
  CLKINVXL U389 ( .A(n60), .Y(n260) );
  CLKINVXL U390 ( .A(n98), .Y(n96) );
  CLKINVXL U391 ( .A(n53), .Y(n259) );
  CLKINVXL U392 ( .A(n80), .Y(n78) );
  CLKINVXL U393 ( .A(n147), .Y(n271) );
  NAND2BXL U394 ( .AN(n136), .B(n137), .Y(n13) );
  NAND2XL U395 ( .A(n270), .B(n142), .Y(n14) );
  CLKINVXL U396 ( .A(n141), .Y(n270) );
  CLKINVXL U397 ( .A(n91), .Y(n263) );
  NAND2XL U398 ( .A(n273), .B(n158), .Y(n17) );
  NAND2XL U399 ( .A(n432), .B(n171), .Y(n19) );
  XOR2X1 U400 ( .A(n180), .B(n424), .Y(SUM[19]) );
  AND2X1 U401 ( .A(n277), .B(n179), .Y(n424) );
  CLKINVXL U402 ( .A(n173), .Y(n276) );
  NAND2XL U403 ( .A(n278), .B(n182), .Y(n22) );
  OAI21XL U404 ( .A0(n195), .A1(n193), .B0(n194), .Y(n192) );
  NAND2XL U405 ( .A(n281), .B(n194), .Y(n25) );
  NAND2XL U406 ( .A(n282), .B(n198), .Y(n26) );
  CLKINVXL U407 ( .A(n193), .Y(n281) );
  NAND2XL U408 ( .A(n431), .B(n203), .Y(n27) );
  CLKINVXL U409 ( .A(n197), .Y(n282) );
  NAND2XL U410 ( .A(n286), .B(n214), .Y(n30) );
  CLKINVXL U411 ( .A(n213), .Y(n286) );
  NAND2XL U412 ( .A(n428), .B(n219), .Y(n31) );
  NAND2XL U413 ( .A(n290), .B(n230), .Y(n34) );
  CLKINVXL U414 ( .A(n229), .Y(n290) );
  NAND2XL U415 ( .A(n430), .B(n239), .Y(n36) );
  INVX1 U416 ( .A(n241), .Y(n293) );
  OR2XL U417 ( .A(B[24]), .B(A[24]), .Y(n429) );
  NAND2XL U418 ( .A(B[8]), .B(A[8]), .Y(n222) );
  OR2XL U419 ( .A(B[7]), .B(A[7]), .Y(n433) );
  NAND2XL U420 ( .A(B[23]), .B(A[23]), .Y(n158) );
  NAND2XL U421 ( .A(B[7]), .B(A[7]), .Y(n227) );
  NAND2XL U422 ( .A(B[11]), .B(A[11]), .Y(n211) );
  NAND2XL U423 ( .A(B[34]), .B(A[34]), .Y(n81) );
  NAND2XL U424 ( .A(B[13]), .B(A[13]), .Y(n203) );
  NAND2XL U425 ( .A(B[30]), .B(A[30]), .Y(n113) );
  NAND2XL U426 ( .A(B[20]), .B(A[20]), .Y(n174) );
  NAND2XL U427 ( .A(B[36]), .B(A[36]), .Y(n63) );
  NAND2XL U428 ( .A(B[17]), .B(A[17]), .Y(n186) );
  NAND2XL U429 ( .A(B[21]), .B(A[21]), .Y(n171) );
  NAND2XL U430 ( .A(B[12]), .B(A[12]), .Y(n206) );
  NAND2XL U431 ( .A(B[22]), .B(A[22]), .Y(n166) );
  NAND2XL U432 ( .A(B[4]), .B(A[4]), .Y(n239) );
  NAND2X1 U433 ( .A(n425), .B(n426), .Y(n1) );
  OR2XL U434 ( .A(n437), .B(A[39]), .Y(n425) );
  NAND2XL U435 ( .A(n437), .B(A[39]), .Y(n426) );
  XNOR2XL U436 ( .A(n36), .B(n240), .Y(SUM[4]) );
  INVX2 U437 ( .A(n438), .Y(n437) );
  INVX2 U438 ( .A(B[38]), .Y(n438) );
  INVX2 U439 ( .A(n83), .Y(n85) );
  NOR2X1 U440 ( .A(n49), .B(n83), .Y(n47) );
  OAI21X1 U441 ( .A0(n84), .A1(n49), .B0(n50), .Y(n48) );
  NAND2X1 U442 ( .A(n67), .B(n51), .Y(n49) );
  INVX2 U443 ( .A(n67), .Y(n69) );
  NAND2X1 U444 ( .A(n85), .B(n67), .Y(n65) );
  OAI21XL U445 ( .A0(n114), .A1(n83), .B0(n84), .Y(n82) );
  INVX2 U446 ( .A(n130), .Y(n132) );
  OAI21XL U447 ( .A0(n114), .A1(n56), .B0(n57), .Y(n55) );
  NOR2X1 U448 ( .A(n69), .B(n60), .Y(n58) );
  XNOR2X1 U449 ( .A(n55), .B(n3), .Y(SUM[37]) );
  NAND2X1 U450 ( .A(n259), .B(n54), .Y(n3) );
  NOR2X1 U451 ( .A(n60), .B(n53), .Y(n51) );
  OAI21X1 U452 ( .A0(n73), .A1(n81), .B0(n74), .Y(n68) );
  NAND2X1 U453 ( .A(n258), .B(n45), .Y(n2) );
  OAI21X1 U454 ( .A0(n199), .A1(n197), .B0(n198), .Y(n196) );
  NAND2X1 U455 ( .A(n130), .B(n118), .Y(n116) );
  OAI21XL U456 ( .A0(n120), .A1(n128), .B0(n121), .Y(n119) );
  OAI21X1 U457 ( .A0(n178), .A1(n182), .B0(n179), .Y(n177) );
  NOR2X1 U458 ( .A(n181), .B(n178), .Y(n176) );
  OAI21X1 U459 ( .A0(n173), .A1(n175), .B0(n174), .Y(n172) );
  NOR2X1 U460 ( .A(n150), .B(n147), .Y(n145) );
  OAI21X1 U461 ( .A0(n187), .A1(n185), .B0(n186), .Y(n184) );
  AOI21X1 U462 ( .A0(n188), .A1(n196), .B0(n189), .Y(n187) );
  OAI21X1 U463 ( .A0(n190), .A1(n194), .B0(n191), .Y(n189) );
  NOR2X1 U464 ( .A(n193), .B(n190), .Y(n188) );
  AOI21X1 U465 ( .A0(n172), .A1(n432), .B0(n169), .Y(n167) );
  INVX2 U466 ( .A(n171), .Y(n169) );
  XNOR2X1 U467 ( .A(n64), .B(n4), .Y(SUM[36]) );
  NAND2X1 U468 ( .A(n260), .B(n63), .Y(n4) );
  XNOR2X1 U469 ( .A(n100), .B(n8), .Y(SUM[32]) );
  OAI21XL U470 ( .A0(n114), .A1(n94), .B0(n95), .Y(n93) );
  NAND2XL U471 ( .A(n103), .B(n96), .Y(n94) );
  XNOR2X1 U472 ( .A(n93), .B(n7), .Y(SUM[33]) );
  NOR2X1 U473 ( .A(n125), .B(n120), .Y(n118) );
  OAI21XL U474 ( .A0(n114), .A1(n112), .B0(n113), .Y(n111) );
  OAI21XL U475 ( .A0(n114), .A1(n76), .B0(n77), .Y(n75) );
  XNOR2X1 U476 ( .A(n82), .B(n6), .Y(SUM[34]) );
  INVX2 U477 ( .A(n203), .Y(n201) );
  OAI21X1 U478 ( .A0(n205), .A1(n207), .B0(n206), .Y(n204) );
  OAI21X1 U479 ( .A0(n142), .A1(n136), .B0(n137), .Y(n131) );
  OAI21X1 U480 ( .A0(n213), .A1(n215), .B0(n214), .Y(n212) );
  AOI21X1 U481 ( .A0(n435), .A1(n212), .B0(n209), .Y(n207) );
  INVX2 U482 ( .A(n211), .Y(n209) );
  INVX2 U483 ( .A(n227), .Y(n225) );
  OAI21X1 U484 ( .A0(n221), .A1(n223), .B0(n222), .Y(n220) );
  OAI21X1 U485 ( .A0(n229), .A1(n231), .B0(n230), .Y(n228) );
  OAI21X1 U486 ( .A0(n233), .A1(n235), .B0(n234), .Y(n232) );
  INVX2 U487 ( .A(n239), .Y(n237) );
  XOR2X1 U488 ( .A(n129), .B(n12), .Y(SUM[28]) );
  OAI21XL U489 ( .A0(n133), .A1(n125), .B0(n128), .Y(n124) );
  NOR2X1 U490 ( .A(n132), .B(n125), .Y(n123) );
  CLKINVXL U491 ( .A(n131), .Y(n133) );
  XOR2X1 U492 ( .A(n122), .B(n11), .Y(SUM[29]) );
  NAND2X1 U493 ( .A(n273), .B(n429), .Y(n150) );
  AOI21X1 U494 ( .A0(n89), .A1(n104), .B0(n90), .Y(n84) );
  OAI21X1 U495 ( .A0(n91), .A1(n99), .B0(n92), .Y(n90) );
  OAI21X1 U496 ( .A0(n109), .A1(n113), .B0(n110), .Y(n104) );
  INVX2 U497 ( .A(n247), .Y(n245) );
  OAI21X1 U498 ( .A0(n241), .A1(n243), .B0(n242), .Y(n240) );
  NOR2X1 U499 ( .A(n91), .B(n98), .Y(n89) );
  OAI2BB1X1 U500 ( .A0N(n436), .A1N(n254), .B0(n253), .Y(n427) );
  XNOR2X1 U501 ( .A(n149), .B(n15), .Y(SUM[25]) );
  NAND2BX1 U502 ( .AN(n73), .B(n74), .Y(n5) );
  CLKINVXL U503 ( .A(n125), .Y(n268) );
  CLKINVXL U504 ( .A(n120), .Y(n267) );
  INVX2 U505 ( .A(n256), .Y(n254) );
  NAND2BX1 U506 ( .AN(n112), .B(n113), .Y(n10) );
  NAND2BX1 U507 ( .AN(n109), .B(n110), .Y(n9) );
  NAND2X1 U508 ( .A(n276), .B(n174), .Y(n20) );
  NAND2BX1 U509 ( .AN(n165), .B(n166), .Y(n18) );
  OAI21XL U510 ( .A0(n183), .A1(n181), .B0(n182), .Y(n180) );
  CLKINVXL U511 ( .A(n181), .Y(n278) );
  XOR2X1 U512 ( .A(n183), .B(n22), .Y(SUM[18]) );
  CLKINVXL U513 ( .A(n178), .Y(n277) );
  NAND2BX1 U514 ( .AN(n185), .B(n186), .Y(n23) );
  XOR2X1 U515 ( .A(n25), .B(n195), .Y(SUM[15]) );
  NAND2BX1 U516 ( .AN(n190), .B(n191), .Y(n24) );
  NAND2BX1 U517 ( .AN(n205), .B(n206), .Y(n28) );
  NAND2X1 U518 ( .A(n435), .B(n211), .Y(n29) );
  NAND2BX1 U519 ( .AN(n221), .B(n222), .Y(n32) );
  XNOR2XL U520 ( .A(n33), .B(n228), .Y(SUM[7]) );
  NAND2X1 U521 ( .A(n433), .B(n227), .Y(n33) );
  XOR2XL U522 ( .A(n34), .B(n231), .Y(SUM[6]) );
  NAND2BX1 U523 ( .AN(n233), .B(n234), .Y(n35) );
  NAND2X1 U524 ( .A(n293), .B(n242), .Y(n37) );
  XNOR2X1 U525 ( .A(n38), .B(n427), .Y(SUM[2]) );
  NAND2X1 U526 ( .A(n434), .B(n247), .Y(n38) );
  NAND2X1 U527 ( .A(n436), .B(n253), .Y(n39) );
  XNOR2X1 U528 ( .A(n43), .B(n1), .Y(SUM[39]) );
  NOR2X1 U529 ( .A(B[34]), .B(A[34]), .Y(n80) );
  NOR2X1 U530 ( .A(B[37]), .B(A[37]), .Y(n53) );
  NOR2X1 U531 ( .A(B[36]), .B(A[36]), .Y(n60) );
  NOR2X1 U532 ( .A(B[14]), .B(A[14]), .Y(n197) );
  NAND2XL U533 ( .A(B[35]), .B(A[35]), .Y(n74) );
  NOR2X1 U534 ( .A(B[26]), .B(A[26]), .Y(n141) );
  NOR2X1 U535 ( .A(B[20]), .B(A[20]), .Y(n173) );
  XNOR2X1 U536 ( .A(n111), .B(n9), .Y(SUM[31]) );
  XNOR2X1 U537 ( .A(n75), .B(n5), .Y(SUM[35]) );
  NOR2X1 U538 ( .A(B[12]), .B(A[12]), .Y(n205) );
  OR2XL U539 ( .A(B[9]), .B(A[9]), .Y(n428) );
  NOR2X1 U540 ( .A(B[5]), .B(A[5]), .Y(n233) );
  NAND2XL U541 ( .A(B[37]), .B(A[37]), .Y(n54) );
  OR2XL U542 ( .A(B[4]), .B(A[4]), .Y(n430) );
  NAND2X1 U543 ( .A(B[18]), .B(A[18]), .Y(n182) );
  OR2X1 U544 ( .A(B[13]), .B(A[13]), .Y(n431) );
  NAND2X1 U545 ( .A(B[26]), .B(A[26]), .Y(n142) );
  NOR2X1 U546 ( .A(n437), .B(A[38]), .Y(n44) );
  NOR2X1 U547 ( .A(B[15]), .B(A[15]), .Y(n193) );
  OR2X1 U548 ( .A(B[21]), .B(A[21]), .Y(n432) );
  NAND2XL U549 ( .A(B[14]), .B(A[14]), .Y(n198) );
  NOR2X1 U550 ( .A(B[25]), .B(A[25]), .Y(n147) );
  NOR2X1 U551 ( .A(B[31]), .B(A[31]), .Y(n109) );
  NOR2X1 U552 ( .A(B[6]), .B(A[6]), .Y(n229) );
  NOR2X1 U553 ( .A(B[17]), .B(A[17]), .Y(n185) );
  NOR2X1 U554 ( .A(B[10]), .B(A[10]), .Y(n213) );
  NAND2XL U555 ( .A(B[27]), .B(A[27]), .Y(n137) );
  NAND2XL U556 ( .A(B[24]), .B(A[24]), .Y(n155) );
  NAND2X1 U557 ( .A(B[15]), .B(A[15]), .Y(n194) );
  XOR2X1 U558 ( .A(n138), .B(n13), .Y(SUM[27]) );
  NAND2XL U559 ( .A(B[19]), .B(A[19]), .Y(n179) );
  NAND2XL U560 ( .A(B[5]), .B(A[5]), .Y(n234) );
  NOR2X1 U561 ( .A(B[23]), .B(A[23]), .Y(n157) );
  NAND2X1 U562 ( .A(B[28]), .B(A[28]), .Y(n128) );
  XOR2X1 U563 ( .A(n114), .B(n10), .Y(SUM[30]) );
  OR2X1 U564 ( .A(B[2]), .B(A[2]), .Y(n434) );
  NOR2X1 U565 ( .A(B[32]), .B(A[32]), .Y(n98) );
  NOR2X1 U566 ( .A(B[3]), .B(A[3]), .Y(n241) );
  NAND2XL U567 ( .A(B[9]), .B(A[9]), .Y(n219) );
  NAND2XL U568 ( .A(B[29]), .B(A[29]), .Y(n121) );
  OR2XL U569 ( .A(B[1]), .B(A[1]), .Y(n436) );
  NAND2XL U570 ( .A(B[6]), .B(A[6]), .Y(n230) );
  NAND2XL U571 ( .A(n437), .B(A[38]), .Y(n45) );
  NAND2XL U572 ( .A(B[16]), .B(A[16]), .Y(n191) );
  NAND2XL U573 ( .A(B[25]), .B(A[25]), .Y(n148) );
  NOR2X1 U574 ( .A(B[8]), .B(A[8]), .Y(n221) );
  NAND2X1 U575 ( .A(B[2]), .B(A[2]), .Y(n247) );
  NAND2XL U576 ( .A(B[10]), .B(A[10]), .Y(n214) );
  NAND2XL U577 ( .A(B[32]), .B(A[32]), .Y(n99) );
  NOR2X1 U578 ( .A(B[33]), .B(A[33]), .Y(n91) );
  NAND2XL U579 ( .A(B[1]), .B(A[1]), .Y(n253) );
  NAND2XL U580 ( .A(B[3]), .B(A[3]), .Y(n242) );
  NAND2XL U581 ( .A(B[31]), .B(A[31]), .Y(n110) );
  NAND2XL U582 ( .A(B[33]), .B(A[33]), .Y(n92) );
  NOR2X1 U583 ( .A(B[22]), .B(A[22]), .Y(n165) );
  XNOR2X1 U584 ( .A(n143), .B(n14), .Y(SUM[26]) );
  XOR2X1 U585 ( .A(n163), .B(n17), .Y(SUM[23]) );
  NAND2X1 U586 ( .A(B[0]), .B(A[0]), .Y(n256) );
  XNOR2X1 U587 ( .A(n192), .B(n24), .Y(SUM[16]) );
  XNOR2XL U588 ( .A(n27), .B(n204), .Y(SUM[13]) );
  XNOR2XL U589 ( .A(n31), .B(n220), .Y(SUM[9]) );
  XNOR2X1 U590 ( .A(n39), .B(n254), .Y(SUM[1]) );
  NAND2BX1 U591 ( .AN(n255), .B(n256), .Y(n40) );
  NOR2X1 U592 ( .A(B[0]), .B(A[0]), .Y(n255) );
  INVX2 U593 ( .A(n40), .Y(SUM[0]) );
  XNOR2XL U594 ( .A(n29), .B(n212), .Y(SUM[11]) );
  XOR2XL U595 ( .A(n37), .B(n243), .Y(SUM[3]) );
  XOR2XL U596 ( .A(n28), .B(n207), .Y(SUM[12]) );
  XNOR2X1 U597 ( .A(n172), .B(n19), .Y(SUM[21]) );
  INVX2 U598 ( .A(n144), .Y(n143) );
  XOR2X1 U599 ( .A(n46), .B(n2), .Y(SUM[38]) );
  XOR2X1 U600 ( .A(n187), .B(n23), .Y(SUM[17]) );
  XOR2XL U601 ( .A(n20), .B(n175), .Y(SUM[20]) );
  OAI21X1 U602 ( .A0(n46), .A1(n44), .B0(n45), .Y(n43) );
  XOR2XL U603 ( .A(n30), .B(n215), .Y(SUM[10]) );
  XOR2XL U604 ( .A(n18), .B(n167), .Y(SUM[22]) );
  XOR2XL U605 ( .A(n26), .B(n199), .Y(SUM[14]) );
  XOR2XL U606 ( .A(n32), .B(n223), .Y(SUM[8]) );
  XOR2XL U607 ( .A(n35), .B(n235), .Y(SUM[5]) );
endmodule


module MMSA_DW01_add_31 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n20, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n63, n64, n65, n66, n67, n68, n69, n70, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n128, n129, n130, n131, n132, n133, n136,
         n137, n138, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n153, n155, n156, n157, n158, n160, n163, n164,
         n165, n166, n167, n169, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n201, n203, n204, n205, n206, n207, n209, n211, n212, n213, n214,
         n215, n217, n219, n220, n221, n222, n223, n225, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n237, n239, n240, n241, n242,
         n243, n245, n247, n253, n254, n255, n256, n258, n259, n260, n263,
         n267, n268, n270, n271, n273, n276, n277, n278, n281, n282, n286,
         n290, n293, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434;

  AOI21X1 U17 ( .A0(n51), .A1(n68), .B0(n52), .Y(n50) );
  AOI21X1 U27 ( .A0(n58), .A1(n86), .B0(n59), .Y(n57) );
  AOI21X1 U39 ( .A0(n86), .A1(n67), .B0(n68), .Y(n66) );
  AOI21X1 U53 ( .A0(n86), .A1(n78), .B0(n79), .Y(n77) );
  AOI21X1 U77 ( .A0(n104), .A1(n96), .B0(n97), .Y(n95) );
  AOI21X1 U108 ( .A0(n131), .A1(n118), .B0(n119), .Y(n117) );
  NOR2X2 U113 ( .A(B[29]), .B(A[29]), .Y(n120) );
  NOR2X2 U123 ( .A(B[28]), .B(A[28]), .Y(n125) );
  AOI21X1 U126 ( .A0(n143), .A1(n130), .B0(n131), .Y(n129) );
  AOI21X1 U138 ( .A0(n143), .A1(n270), .B0(n140), .Y(n138) );
  AOI21X1 U157 ( .A0(n427), .A1(n160), .B0(n153), .Y(n151) );
  OAI21XL U340 ( .A0(n190), .A1(n194), .B0(n191), .Y(n189) );
  OAI21X2 U341 ( .A0(n173), .A1(n175), .B0(n174), .Y(n172) );
  OAI21X2 U342 ( .A0(n187), .A1(n185), .B0(n186), .Y(n184) );
  OAI21X2 U343 ( .A0(n116), .A1(n144), .B0(n117), .Y(n115) );
  NOR2XL U344 ( .A(B[35]), .B(A[35]), .Y(n73) );
  NOR2X1 U345 ( .A(n91), .B(n98), .Y(n89) );
  AOI21X1 U346 ( .A0(n145), .A1(n164), .B0(n146), .Y(n144) );
  OAI21X2 U347 ( .A0(n165), .A1(n167), .B0(n166), .Y(n164) );
  NOR2X1 U348 ( .A(B[19]), .B(A[19]), .Y(n178) );
  NOR2X1 U349 ( .A(B[18]), .B(A[18]), .Y(n181) );
  NAND2X1 U350 ( .A(n130), .B(n118), .Y(n116) );
  AOI21X1 U351 ( .A0(n89), .A1(n104), .B0(n90), .Y(n84) );
  NOR2X1 U352 ( .A(n80), .B(n73), .Y(n67) );
  OAI21X1 U353 ( .A0(n109), .A1(n113), .B0(n110), .Y(n104) );
  NOR2X1 U354 ( .A(n112), .B(n109), .Y(n103) );
  NOR2X1 U355 ( .A(B[27]), .B(A[27]), .Y(n136) );
  NOR2X1 U356 ( .A(B[30]), .B(A[30]), .Y(n112) );
  INVX2 U357 ( .A(n115), .Y(n114) );
  OAI21X1 U358 ( .A0(n91), .A1(n99), .B0(n92), .Y(n90) );
  AOI21X1 U359 ( .A0(n123), .A1(n143), .B0(n124), .Y(n122) );
  OAI21X1 U360 ( .A0(n114), .A1(n65), .B0(n66), .Y(n64) );
  NAND2XL U361 ( .A(n85), .B(n67), .Y(n65) );
  OAI21XL U362 ( .A0(n114), .A1(n101), .B0(n102), .Y(n100) );
  CLKINVX2 U363 ( .A(n84), .Y(n86) );
  OAI21X1 U364 ( .A0(n70), .A1(n60), .B0(n63), .Y(n59) );
  CLKINVXL U365 ( .A(n103), .Y(n101) );
  OAI21XL U366 ( .A0(n163), .A1(n150), .B0(n151), .Y(n149) );
  NAND2X1 U367 ( .A(n89), .B(n103), .Y(n83) );
  CLKINVXL U368 ( .A(n130), .Y(n132) );
  CLKINVXL U369 ( .A(n196), .Y(n195) );
  OAI21X1 U370 ( .A0(n151), .A1(n147), .B0(n148), .Y(n146) );
  NAND2XL U371 ( .A(n267), .B(n121), .Y(n11) );
  CLKINVX2 U372 ( .A(n99), .Y(n97) );
  OAI21XL U373 ( .A0(n114), .A1(n94), .B0(n95), .Y(n93) );
  OAI21XL U374 ( .A0(n114), .A1(n56), .B0(n57), .Y(n55) );
  NAND2XL U375 ( .A(n78), .B(n81), .Y(n6) );
  CLKINVXL U376 ( .A(n81), .Y(n79) );
  NAND2XL U377 ( .A(n85), .B(n78), .Y(n76) );
  OAI21X1 U378 ( .A0(n142), .A1(n136), .B0(n137), .Y(n131) );
  NAND2XL U379 ( .A(n271), .B(n148), .Y(n15) );
  CLKINVX2 U380 ( .A(n157), .Y(n273) );
  INVX1 U381 ( .A(n68), .Y(n70) );
  OAI21XL U382 ( .A0(n53), .A1(n63), .B0(n54), .Y(n52) );
  OAI21XL U383 ( .A0(n163), .A1(n157), .B0(n158), .Y(n156) );
  INVX1 U384 ( .A(n232), .Y(n231) );
  CLKINVXL U385 ( .A(n60), .Y(n260) );
  CLKINVXL U386 ( .A(n53), .Y(n259) );
  CLKINVXL U387 ( .A(n80), .Y(n78) );
  CLKINVXL U388 ( .A(n98), .Y(n96) );
  CLKINVXL U389 ( .A(n147), .Y(n271) );
  NAND2XL U390 ( .A(n270), .B(n142), .Y(n14) );
  CLKINVXL U391 ( .A(n141), .Y(n270) );
  CLKINVXL U392 ( .A(n91), .Y(n263) );
  NAND2BXL U393 ( .AN(n112), .B(n113), .Y(n10) );
  XOR2X1 U394 ( .A(n172), .B(n423), .Y(SUM[21]) );
  AND2X1 U395 ( .A(n432), .B(n171), .Y(n423) );
  NAND2XL U396 ( .A(n276), .B(n174), .Y(n20) );
  XOR2X1 U397 ( .A(n180), .B(n424), .Y(SUM[19]) );
  AND2X1 U398 ( .A(n277), .B(n179), .Y(n424) );
  CLKINVXL U399 ( .A(n173), .Y(n276) );
  OAI21XL U400 ( .A0(n195), .A1(n193), .B0(n194), .Y(n192) );
  NAND2XL U401 ( .A(n282), .B(n198), .Y(n26) );
  CLKINVXL U402 ( .A(n193), .Y(n281) );
  CLKINVXL U403 ( .A(n197), .Y(n282) );
  NAND2XL U404 ( .A(n286), .B(n214), .Y(n30) );
  CLKINVXL U405 ( .A(n213), .Y(n286) );
  NAND2XL U406 ( .A(n430), .B(n227), .Y(n33) );
  NAND2XL U407 ( .A(n290), .B(n230), .Y(n34) );
  CLKINVXL U408 ( .A(n229), .Y(n290) );
  OR2XL U409 ( .A(B[24]), .B(A[24]), .Y(n427) );
  NAND2XL U410 ( .A(B[24]), .B(A[24]), .Y(n155) );
  NAND2XL U411 ( .A(B[23]), .B(A[23]), .Y(n158) );
  NAND2XL U412 ( .A(B[8]), .B(A[8]), .Y(n222) );
  OR2XL U413 ( .A(B[11]), .B(A[11]), .Y(n431) );
  OR2XL U414 ( .A(B[7]), .B(A[7]), .Y(n430) );
  NAND2XL U415 ( .A(B[11]), .B(A[11]), .Y(n211) );
  OR2XL U416 ( .A(B[13]), .B(A[13]), .Y(n433) );
  NAND2XL U417 ( .A(B[18]), .B(A[18]), .Y(n182) );
  OR2XL U418 ( .A(B[21]), .B(A[21]), .Y(n432) );
  NAND2XL U419 ( .A(B[28]), .B(A[28]), .Y(n128) );
  NAND2XL U420 ( .A(B[15]), .B(A[15]), .Y(n194) );
  NAND2XL U421 ( .A(B[13]), .B(A[13]), .Y(n203) );
  NAND2XL U422 ( .A(B[21]), .B(A[21]), .Y(n171) );
  NAND2XL U423 ( .A(B[22]), .B(A[22]), .Y(n166) );
  OR2XL U424 ( .A(B[4]), .B(A[4]), .Y(n426) );
  NAND2XL U425 ( .A(B[4]), .B(A[4]), .Y(n239) );
  NAND2BX1 U426 ( .AN(n41), .B(n42), .Y(n1) );
  INVX2 U427 ( .A(n83), .Y(n85) );
  AOI21X1 U428 ( .A0(n115), .A1(n47), .B0(n48), .Y(n46) );
  OAI21X1 U429 ( .A0(n84), .A1(n49), .B0(n50), .Y(n48) );
  NAND2X1 U430 ( .A(n67), .B(n51), .Y(n49) );
  INVX2 U431 ( .A(n67), .Y(n69) );
  INVX2 U432 ( .A(n104), .Y(n102) );
  OAI21XL U433 ( .A0(n114), .A1(n83), .B0(n84), .Y(n82) );
  INVX2 U434 ( .A(n144), .Y(n143) );
  INVX2 U435 ( .A(n164), .Y(n163) );
  INVX2 U436 ( .A(n184), .Y(n183) );
  OAI21X1 U437 ( .A0(n46), .A1(n44), .B0(n45), .Y(n43) );
  XNOR2X1 U438 ( .A(n55), .B(n3), .Y(SUM[37]) );
  NAND2X1 U439 ( .A(n259), .B(n54), .Y(n3) );
  NAND2X1 U440 ( .A(n58), .B(n85), .Y(n56) );
  NOR2X1 U441 ( .A(n69), .B(n60), .Y(n58) );
  XOR2X1 U442 ( .A(n46), .B(n2), .Y(SUM[38]) );
  NAND2X1 U443 ( .A(n258), .B(n45), .Y(n2) );
  NOR2X1 U444 ( .A(n60), .B(n53), .Y(n51) );
  XNOR2X1 U445 ( .A(n64), .B(n4), .Y(SUM[36]) );
  NAND2X1 U446 ( .A(n260), .B(n63), .Y(n4) );
  XNOR2X1 U447 ( .A(n100), .B(n8), .Y(SUM[32]) );
  NAND2X1 U448 ( .A(n96), .B(n99), .Y(n8) );
  XNOR2X1 U449 ( .A(n93), .B(n7), .Y(SUM[33]) );
  NAND2X1 U450 ( .A(n263), .B(n92), .Y(n7) );
  NOR2X1 U451 ( .A(n141), .B(n136), .Y(n130) );
  OAI21XL U452 ( .A0(n120), .A1(n128), .B0(n121), .Y(n119) );
  NAND2XL U453 ( .A(n103), .B(n96), .Y(n94) );
  NOR2X1 U454 ( .A(n150), .B(n147), .Y(n145) );
  AOI21X1 U455 ( .A0(n172), .A1(n432), .B0(n169), .Y(n167) );
  INVX2 U456 ( .A(n171), .Y(n169) );
  OAI21X1 U457 ( .A0(n205), .A1(n207), .B0(n206), .Y(n204) );
  OAI21X1 U458 ( .A0(n229), .A1(n231), .B0(n230), .Y(n228) );
  AOI21X1 U459 ( .A0(n204), .A1(n433), .B0(n201), .Y(n199) );
  INVX2 U460 ( .A(n203), .Y(n201) );
  AOI21X1 U461 ( .A0(n426), .A1(n240), .B0(n237), .Y(n235) );
  INVX2 U462 ( .A(n239), .Y(n237) );
  AOI21X1 U463 ( .A0(n176), .A1(n184), .B0(n177), .Y(n175) );
  OAI21X1 U464 ( .A0(n178), .A1(n182), .B0(n179), .Y(n177) );
  NOR2X1 U465 ( .A(n181), .B(n178), .Y(n176) );
  AOI21X1 U466 ( .A0(n228), .A1(n430), .B0(n225), .Y(n223) );
  INVX2 U467 ( .A(n227), .Y(n225) );
  OAI21X1 U468 ( .A0(n221), .A1(n223), .B0(n222), .Y(n220) );
  OAI21X1 U469 ( .A0(n199), .A1(n197), .B0(n198), .Y(n196) );
  AOI21X1 U470 ( .A0(n431), .A1(n212), .B0(n209), .Y(n207) );
  INVX2 U471 ( .A(n211), .Y(n209) );
  AOI21X1 U472 ( .A0(n188), .A1(n196), .B0(n189), .Y(n187) );
  NOR2X1 U473 ( .A(n193), .B(n190), .Y(n188) );
  OAI21X1 U474 ( .A0(n213), .A1(n215), .B0(n214), .Y(n212) );
  AOI21X1 U475 ( .A0(n220), .A1(n434), .B0(n217), .Y(n215) );
  INVX2 U476 ( .A(n219), .Y(n217) );
  OAI21X1 U477 ( .A0(n233), .A1(n235), .B0(n234), .Y(n232) );
  NOR2X1 U478 ( .A(n125), .B(n120), .Y(n118) );
  OAI21X1 U479 ( .A0(n73), .A1(n81), .B0(n74), .Y(n68) );
  XNOR2X1 U480 ( .A(n82), .B(n6), .Y(SUM[34]) );
  OAI21XL U481 ( .A0(n114), .A1(n112), .B0(n113), .Y(n111) );
  OAI21XL U482 ( .A0(n114), .A1(n76), .B0(n77), .Y(n75) );
  NAND2X1 U483 ( .A(n273), .B(n427), .Y(n150) );
  XOR2X1 U484 ( .A(n129), .B(n12), .Y(SUM[28]) );
  NAND2X1 U485 ( .A(n268), .B(n128), .Y(n12) );
  INVX2 U486 ( .A(n155), .Y(n153) );
  INVX2 U487 ( .A(n158), .Y(n160) );
  AOI21X1 U488 ( .A0(n428), .A1(n425), .B0(n245), .Y(n243) );
  INVX2 U489 ( .A(n247), .Y(n245) );
  OAI21X1 U490 ( .A0(n241), .A1(n243), .B0(n242), .Y(n240) );
  OAI2BB1X1 U491 ( .A0N(n429), .A1N(n254), .B0(n253), .Y(n425) );
  INVX2 U492 ( .A(n142), .Y(n140) );
  OAI21XL U493 ( .A0(n133), .A1(n125), .B0(n128), .Y(n124) );
  NOR2X1 U494 ( .A(n132), .B(n125), .Y(n123) );
  CLKINVXL U495 ( .A(n131), .Y(n133) );
  XOR2X1 U496 ( .A(n122), .B(n11), .Y(SUM[29]) );
  INVX2 U497 ( .A(n44), .Y(n258) );
  XNOR2X1 U498 ( .A(n156), .B(n16), .Y(SUM[24]) );
  NAND2X1 U499 ( .A(n427), .B(n155), .Y(n16) );
  XNOR2X1 U500 ( .A(n149), .B(n15), .Y(SUM[25]) );
  NAND2BX1 U501 ( .AN(n73), .B(n74), .Y(n5) );
  CLKINVXL U502 ( .A(n125), .Y(n268) );
  CLKINVXL U503 ( .A(n120), .Y(n267) );
  NAND2BX1 U504 ( .AN(n136), .B(n137), .Y(n13) );
  INVX2 U505 ( .A(n256), .Y(n254) );
  NAND2BX1 U506 ( .AN(n109), .B(n110), .Y(n9) );
  NAND2XL U507 ( .A(n273), .B(n158), .Y(n17) );
  OAI21XL U508 ( .A0(n183), .A1(n181), .B0(n182), .Y(n180) );
  XOR2XL U509 ( .A(n20), .B(n175), .Y(SUM[20]) );
  XOR2X1 U510 ( .A(n183), .B(n22), .Y(SUM[18]) );
  NAND2X1 U511 ( .A(n278), .B(n182), .Y(n22) );
  NAND2BX1 U512 ( .AN(n165), .B(n166), .Y(n18) );
  CLKINVXL U513 ( .A(n181), .Y(n278) );
  CLKINVXL U514 ( .A(n178), .Y(n277) );
  NAND2BX1 U515 ( .AN(n185), .B(n186), .Y(n23) );
  XOR2X1 U516 ( .A(n25), .B(n195), .Y(SUM[15]) );
  NAND2X1 U517 ( .A(n281), .B(n194), .Y(n25) );
  NAND2BX1 U518 ( .AN(n190), .B(n191), .Y(n24) );
  XOR2XL U519 ( .A(n26), .B(n199), .Y(SUM[14]) );
  NAND2X1 U520 ( .A(n433), .B(n203), .Y(n27) );
  NAND2BX1 U521 ( .AN(n205), .B(n206), .Y(n28) );
  NAND2X1 U522 ( .A(n431), .B(n211), .Y(n29) );
  NAND2XL U523 ( .A(n434), .B(n219), .Y(n31) );
  NAND2BX1 U524 ( .AN(n221), .B(n222), .Y(n32) );
  XNOR2XL U525 ( .A(n33), .B(n228), .Y(SUM[7]) );
  XOR2XL U526 ( .A(n34), .B(n231), .Y(SUM[6]) );
  NAND2BX1 U527 ( .AN(n233), .B(n234), .Y(n35) );
  NAND2X1 U528 ( .A(n426), .B(n239), .Y(n36) );
  XOR2XL U529 ( .A(n37), .B(n243), .Y(SUM[3]) );
  NAND2X1 U530 ( .A(n293), .B(n242), .Y(n37) );
  INVX2 U531 ( .A(n241), .Y(n293) );
  XNOR2XL U532 ( .A(n38), .B(n425), .Y(SUM[2]) );
  NAND2X1 U533 ( .A(n428), .B(n247), .Y(n38) );
  NAND2X1 U534 ( .A(n429), .B(n253), .Y(n39) );
  XNOR2X1 U535 ( .A(n43), .B(n1), .Y(SUM[39]) );
  NOR2X1 U536 ( .A(B[34]), .B(A[34]), .Y(n80) );
  NOR2X1 U537 ( .A(B[37]), .B(A[37]), .Y(n53) );
  NOR2X1 U538 ( .A(B[36]), .B(A[36]), .Y(n60) );
  NOR2X1 U539 ( .A(B[25]), .B(A[25]), .Y(n147) );
  NOR2X1 U540 ( .A(B[5]), .B(A[5]), .Y(n233) );
  XNOR2X1 U541 ( .A(n111), .B(n9), .Y(SUM[31]) );
  XNOR2X1 U542 ( .A(n75), .B(n5), .Y(SUM[35]) );
  NOR2X1 U543 ( .A(B[23]), .B(A[23]), .Y(n157) );
  NAND2XL U544 ( .A(B[34]), .B(A[34]), .Y(n81) );
  NOR2X1 U545 ( .A(B[26]), .B(A[26]), .Y(n141) );
  NOR2X1 U546 ( .A(B[6]), .B(A[6]), .Y(n229) );
  NOR2X1 U547 ( .A(B[12]), .B(A[12]), .Y(n205) );
  NOR2X1 U548 ( .A(B[20]), .B(A[20]), .Y(n173) );
  NOR2X1 U549 ( .A(B[14]), .B(A[14]), .Y(n197) );
  XOR2X1 U550 ( .A(n114), .B(n10), .Y(SUM[30]) );
  OR2X1 U551 ( .A(B[2]), .B(A[2]), .Y(n428) );
  NAND2X1 U552 ( .A(B[26]), .B(A[26]), .Y(n142) );
  OR2XL U553 ( .A(B[1]), .B(A[1]), .Y(n429) );
  NAND2XL U554 ( .A(B[5]), .B(A[5]), .Y(n234) );
  NOR2X1 U555 ( .A(B[16]), .B(A[16]), .Y(n190) );
  NOR2X1 U556 ( .A(B[31]), .B(A[31]), .Y(n109) );
  NAND2XL U557 ( .A(B[35]), .B(A[35]), .Y(n74) );
  NOR2X1 U558 ( .A(B[3]), .B(A[3]), .Y(n241) );
  XOR2X1 U559 ( .A(n138), .B(n13), .Y(SUM[27]) );
  NAND2XL U560 ( .A(B[36]), .B(A[36]), .Y(n63) );
  NOR2X1 U561 ( .A(B[10]), .B(A[10]), .Y(n213) );
  NAND2XL U562 ( .A(B[27]), .B(A[27]), .Y(n137) );
  NOR2X1 U563 ( .A(B[15]), .B(A[15]), .Y(n193) );
  OR2XL U564 ( .A(B[9]), .B(A[9]), .Y(n434) );
  NAND2XL U565 ( .A(B[20]), .B(A[20]), .Y(n174) );
  NAND2XL U566 ( .A(B[37]), .B(A[37]), .Y(n54) );
  NOR2X1 U567 ( .A(B[17]), .B(A[17]), .Y(n185) );
  NOR2X1 U568 ( .A(B[33]), .B(A[33]), .Y(n91) );
  NAND2X1 U569 ( .A(B[2]), .B(A[2]), .Y(n247) );
  NAND2XL U570 ( .A(B[19]), .B(A[19]), .Y(n179) );
  NAND2XL U571 ( .A(B[6]), .B(A[6]), .Y(n230) );
  NAND2XL U572 ( .A(B[12]), .B(A[12]), .Y(n206) );
  NOR2X1 U573 ( .A(B[32]), .B(A[32]), .Y(n98) );
  NAND2XL U574 ( .A(B[14]), .B(A[14]), .Y(n198) );
  NOR2X1 U575 ( .A(B[38]), .B(A[38]), .Y(n44) );
  NAND2XL U576 ( .A(B[7]), .B(A[7]), .Y(n227) );
  NAND2X1 U577 ( .A(B[30]), .B(A[30]), .Y(n113) );
  NAND2XL U578 ( .A(B[29]), .B(A[29]), .Y(n121) );
  NAND2XL U579 ( .A(B[10]), .B(A[10]), .Y(n214) );
  NAND2XL U580 ( .A(B[3]), .B(A[3]), .Y(n242) );
  NAND2XL U581 ( .A(B[1]), .B(A[1]), .Y(n253) );
  NOR2X1 U582 ( .A(B[8]), .B(A[8]), .Y(n221) );
  NAND2X1 U583 ( .A(B[38]), .B(A[39]), .Y(n42) );
  NOR2X1 U584 ( .A(B[38]), .B(A[39]), .Y(n41) );
  NAND2X1 U585 ( .A(B[38]), .B(A[38]), .Y(n45) );
  NAND2XL U586 ( .A(B[25]), .B(A[25]), .Y(n148) );
  NAND2XL U587 ( .A(B[16]), .B(A[16]), .Y(n191) );
  NAND2XL U588 ( .A(B[17]), .B(A[17]), .Y(n186) );
  NAND2XL U589 ( .A(B[32]), .B(A[32]), .Y(n99) );
  NAND2XL U590 ( .A(B[31]), .B(A[31]), .Y(n110) );
  XNOR2X1 U591 ( .A(n143), .B(n14), .Y(SUM[26]) );
  NAND2XL U592 ( .A(B[33]), .B(A[33]), .Y(n92) );
  XOR2X1 U593 ( .A(n163), .B(n17), .Y(SUM[23]) );
  NOR2X1 U594 ( .A(B[22]), .B(A[22]), .Y(n165) );
  XOR2XL U595 ( .A(n18), .B(n167), .Y(SUM[22]) );
  NAND2X1 U596 ( .A(B[0]), .B(A[0]), .Y(n256) );
  XNOR2X1 U597 ( .A(n192), .B(n24), .Y(SUM[16]) );
  XOR2X1 U598 ( .A(n187), .B(n23), .Y(SUM[17]) );
  XNOR2XL U599 ( .A(n27), .B(n204), .Y(SUM[13]) );
  XOR2XL U600 ( .A(n28), .B(n207), .Y(SUM[12]) );
  XNOR2XL U601 ( .A(n31), .B(n220), .Y(SUM[9]) );
  XOR2XL U602 ( .A(n32), .B(n223), .Y(SUM[8]) );
  XOR2XL U603 ( .A(n35), .B(n235), .Y(SUM[5]) );
  XNOR2XL U604 ( .A(n36), .B(n240), .Y(SUM[4]) );
  XNOR2X1 U605 ( .A(n39), .B(n254), .Y(SUM[1]) );
  INVX2 U606 ( .A(n40), .Y(SUM[0]) );
  NAND2BX1 U607 ( .AN(n255), .B(n256), .Y(n40) );
  NOR2X1 U608 ( .A(B[0]), .B(A[0]), .Y(n255) );
  XNOR2XL U609 ( .A(n29), .B(n212), .Y(SUM[11]) );
  XOR2XL U610 ( .A(n30), .B(n215), .Y(SUM[10]) );
  NAND2XL U611 ( .A(B[9]), .B(A[9]), .Y(n219) );
  NOR2X1 U612 ( .A(n49), .B(n83), .Y(n47) );
endmodule


module MMSA_DW01_add_30 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n63, n64, n65, n66, n67, n68, n69, n70, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n128, n129, n130, n131, n132, n133, n136,
         n137, n138, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n153, n155, n156, n157, n158, n160, n163, n164,
         n165, n166, n167, n169, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n201, n203, n204, n205, n206, n207, n209, n211, n212, n213, n214,
         n215, n217, n219, n220, n221, n222, n223, n225, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n237, n239, n240, n241, n242,
         n243, n245, n247, n253, n254, n255, n256, n258, n259, n260, n263,
         n267, n268, n270, n271, n273, n276, n277, n278, n281, n282, n286,
         n290, n293, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434;

  AOI21X1 U17 ( .A0(n51), .A1(n68), .B0(n52), .Y(n50) );
  AOI21X1 U27 ( .A0(n58), .A1(n86), .B0(n59), .Y(n57) );
  AOI21X1 U39 ( .A0(n86), .A1(n67), .B0(n68), .Y(n66) );
  AOI21X1 U53 ( .A0(n86), .A1(n78), .B0(n79), .Y(n77) );
  AOI21X1 U77 ( .A0(n104), .A1(n96), .B0(n97), .Y(n95) );
  OAI21X4 U106 ( .A0(n116), .A1(n144), .B0(n117), .Y(n115) );
  AOI21X1 U108 ( .A0(n131), .A1(n118), .B0(n119), .Y(n117) );
  NOR2X2 U113 ( .A(B[29]), .B(A[29]), .Y(n120) );
  AOI21X1 U116 ( .A0(n123), .A1(n143), .B0(n124), .Y(n122) );
  NOR2X2 U123 ( .A(B[28]), .B(A[28]), .Y(n125) );
  AOI21X1 U126 ( .A0(n143), .A1(n130), .B0(n131), .Y(n129) );
  AOI21X1 U138 ( .A0(n143), .A1(n270), .B0(n140), .Y(n138) );
  AOI21X1 U157 ( .A0(n428), .A1(n160), .B0(n153), .Y(n151) );
  AOI21X1 U252 ( .A0(n427), .A1(n212), .B0(n209), .Y(n207) );
  NOR2XL U340 ( .A(B[35]), .B(A[35]), .Y(n73) );
  NOR2X1 U341 ( .A(B[19]), .B(A[19]), .Y(n178) );
  NOR2X1 U342 ( .A(B[18]), .B(A[18]), .Y(n181) );
  NOR2X1 U343 ( .A(B[34]), .B(A[34]), .Y(n80) );
  NOR2X1 U344 ( .A(n60), .B(n53), .Y(n51) );
  AOI21X1 U345 ( .A0(n89), .A1(n104), .B0(n90), .Y(n84) );
  NAND2X1 U346 ( .A(n130), .B(n118), .Y(n116) );
  OAI21X1 U347 ( .A0(n73), .A1(n81), .B0(n74), .Y(n68) );
  NOR2X1 U348 ( .A(n80), .B(n73), .Y(n67) );
  OAI21X1 U349 ( .A0(n109), .A1(n113), .B0(n110), .Y(n104) );
  NOR2X1 U350 ( .A(n112), .B(n109), .Y(n103) );
  NOR2X1 U351 ( .A(B[36]), .B(A[36]), .Y(n60) );
  NOR2X1 U352 ( .A(B[27]), .B(A[27]), .Y(n136) );
  NOR2X1 U353 ( .A(B[30]), .B(A[30]), .Y(n112) );
  OAI21X1 U354 ( .A0(n165), .A1(n167), .B0(n166), .Y(n164) );
  INVXL U355 ( .A(n155), .Y(n153) );
  NAND2XL U356 ( .A(B[18]), .B(A[18]), .Y(n182) );
  OR2XL U357 ( .A(B[13]), .B(A[13]), .Y(n432) );
  OR2XL U358 ( .A(B[11]), .B(A[11]), .Y(n427) );
  OR2XL U359 ( .A(B[21]), .B(A[21]), .Y(n429) );
  OAI21X1 U360 ( .A0(n114), .A1(n65), .B0(n66), .Y(n64) );
  NAND2XL U361 ( .A(n85), .B(n67), .Y(n65) );
  INVX4 U362 ( .A(n115), .Y(n114) );
  OAI21XL U363 ( .A0(n114), .A1(n101), .B0(n102), .Y(n100) );
  CLKINVX2 U364 ( .A(n84), .Y(n86) );
  CLKINVXL U365 ( .A(n144), .Y(n143) );
  CLKINVX1 U366 ( .A(n158), .Y(n160) );
  CLKINVXL U367 ( .A(n103), .Y(n101) );
  OAI21XL U368 ( .A0(n163), .A1(n150), .B0(n151), .Y(n149) );
  NAND2X1 U369 ( .A(n67), .B(n51), .Y(n49) );
  NAND2X1 U370 ( .A(n89), .B(n103), .Y(n83) );
  INVX1 U371 ( .A(n67), .Y(n69) );
  CLKINVXL U372 ( .A(n130), .Y(n132) );
  CLKINVXL U373 ( .A(n184), .Y(n183) );
  CLKINVXL U374 ( .A(n196), .Y(n195) );
  NAND2XL U375 ( .A(n96), .B(n99), .Y(n8) );
  CLKINVXL U376 ( .A(n99), .Y(n97) );
  OAI21XL U377 ( .A0(n114), .A1(n94), .B0(n95), .Y(n93) );
  NAND2XL U378 ( .A(n263), .B(n92), .Y(n7) );
  OAI21XL U379 ( .A0(n114), .A1(n56), .B0(n57), .Y(n55) );
  NAND2XL U380 ( .A(n267), .B(n121), .Y(n11) );
  NAND2XL U381 ( .A(n78), .B(n81), .Y(n6) );
  NAND2XL U382 ( .A(n85), .B(n78), .Y(n76) );
  OAI21X1 U383 ( .A0(n142), .A1(n136), .B0(n137), .Y(n131) );
  NAND2XL U384 ( .A(n271), .B(n148), .Y(n15) );
  OAI21X1 U385 ( .A0(n70), .A1(n60), .B0(n63), .Y(n59) );
  INVX1 U386 ( .A(n68), .Y(n70) );
  CLKINVX2 U387 ( .A(n157), .Y(n273) );
  OAI21XL U388 ( .A0(n53), .A1(n63), .B0(n54), .Y(n52) );
  XOR2X1 U389 ( .A(n156), .B(n423), .Y(SUM[24]) );
  AND2X1 U390 ( .A(n428), .B(n155), .Y(n423) );
  OAI21XL U391 ( .A0(n163), .A1(n157), .B0(n158), .Y(n156) );
  INVX1 U392 ( .A(n232), .Y(n231) );
  CLKINVXL U393 ( .A(n53), .Y(n259) );
  CLKINVX1 U394 ( .A(n239), .Y(n237) );
  CLKINVXL U395 ( .A(n98), .Y(n96) );
  CLKINVXL U396 ( .A(n147), .Y(n271) );
  NAND2XL U397 ( .A(n270), .B(n142), .Y(n14) );
  CLKINVXL U398 ( .A(n141), .Y(n270) );
  CLKINVXL U399 ( .A(n91), .Y(n263) );
  NAND2BXL U400 ( .AN(n112), .B(n113), .Y(n10) );
  NAND2XL U401 ( .A(n276), .B(n174), .Y(n20) );
  XOR2X1 U402 ( .A(n180), .B(n424), .Y(SUM[19]) );
  AND2X1 U403 ( .A(n277), .B(n179), .Y(n424) );
  CLKINVXL U404 ( .A(n173), .Y(n276) );
  OAI21XL U405 ( .A0(n195), .A1(n193), .B0(n194), .Y(n192) );
  NAND2XL U406 ( .A(n282), .B(n198), .Y(n26) );
  CLKINVXL U407 ( .A(n193), .Y(n281) );
  CLKINVXL U408 ( .A(n197), .Y(n282) );
  NAND2XL U409 ( .A(n286), .B(n214), .Y(n30) );
  CLKINVXL U410 ( .A(n213), .Y(n286) );
  NAND2XL U411 ( .A(n431), .B(n219), .Y(n31) );
  NAND2XL U412 ( .A(n290), .B(n230), .Y(n34) );
  CLKINVXL U413 ( .A(n229), .Y(n290) );
  NAND2XL U414 ( .A(n426), .B(n239), .Y(n36) );
  OR2XL U415 ( .A(B[24]), .B(A[24]), .Y(n428) );
  NAND2XL U416 ( .A(B[23]), .B(A[23]), .Y(n158) );
  NAND2XL U417 ( .A(B[8]), .B(A[8]), .Y(n222) );
  NAND2XL U418 ( .A(B[34]), .B(A[34]), .Y(n81) );
  OR2XL U419 ( .A(B[7]), .B(A[7]), .Y(n430) );
  NAND2XL U420 ( .A(B[7]), .B(A[7]), .Y(n227) );
  NAND2XL U421 ( .A(B[11]), .B(A[11]), .Y(n211) );
  NAND2XL U422 ( .A(B[28]), .B(A[28]), .Y(n128) );
  NAND2XL U423 ( .A(B[13]), .B(A[13]), .Y(n203) );
  NAND2XL U424 ( .A(B[15]), .B(A[15]), .Y(n194) );
  NAND2XL U425 ( .A(B[17]), .B(A[17]), .Y(n186) );
  NAND2XL U426 ( .A(B[21]), .B(A[21]), .Y(n171) );
  OR2XL U427 ( .A(B[4]), .B(A[4]), .Y(n426) );
  NAND2XL U428 ( .A(B[22]), .B(A[22]), .Y(n166) );
  NAND2BX1 U429 ( .AN(n41), .B(n42), .Y(n1) );
  INVX2 U430 ( .A(n83), .Y(n85) );
  AOI21X1 U431 ( .A0(n115), .A1(n47), .B0(n48), .Y(n46) );
  OAI21X1 U432 ( .A0(n84), .A1(n49), .B0(n50), .Y(n48) );
  INVX2 U433 ( .A(n104), .Y(n102) );
  OAI21XL U434 ( .A0(n114), .A1(n83), .B0(n84), .Y(n82) );
  INVX2 U435 ( .A(n164), .Y(n163) );
  OAI21X1 U436 ( .A0(n46), .A1(n44), .B0(n45), .Y(n43) );
  XNOR2X1 U437 ( .A(n55), .B(n3), .Y(SUM[37]) );
  NAND2X1 U438 ( .A(n259), .B(n54), .Y(n3) );
  NAND2X1 U439 ( .A(n58), .B(n85), .Y(n56) );
  NOR2X1 U440 ( .A(n69), .B(n60), .Y(n58) );
  XOR2X1 U441 ( .A(n46), .B(n2), .Y(SUM[38]) );
  NAND2X1 U442 ( .A(n258), .B(n45), .Y(n2) );
  XNOR2X1 U443 ( .A(n64), .B(n4), .Y(SUM[36]) );
  NAND2X1 U444 ( .A(n260), .B(n63), .Y(n4) );
  NOR2X1 U445 ( .A(n141), .B(n136), .Y(n130) );
  OAI21XL U446 ( .A0(n120), .A1(n128), .B0(n121), .Y(n119) );
  XNOR2X1 U447 ( .A(n100), .B(n8), .Y(SUM[32]) );
  XNOR2X1 U448 ( .A(n93), .B(n7), .Y(SUM[33]) );
  NAND2XL U449 ( .A(n103), .B(n96), .Y(n94) );
  NOR2X1 U450 ( .A(n125), .B(n120), .Y(n118) );
  AOI21X1 U451 ( .A0(n176), .A1(n184), .B0(n177), .Y(n175) );
  OAI21X1 U452 ( .A0(n178), .A1(n182), .B0(n179), .Y(n177) );
  NOR2X1 U453 ( .A(n181), .B(n178), .Y(n176) );
  AOI21X1 U454 ( .A0(n172), .A1(n429), .B0(n169), .Y(n167) );
  INVX2 U455 ( .A(n171), .Y(n169) );
  AOI21X2 U456 ( .A0(n145), .A1(n164), .B0(n146), .Y(n144) );
  OAI21X1 U457 ( .A0(n151), .A1(n147), .B0(n148), .Y(n146) );
  OAI21X1 U458 ( .A0(n173), .A1(n175), .B0(n174), .Y(n172) );
  XNOR2X1 U459 ( .A(n82), .B(n6), .Y(SUM[34]) );
  OAI21XL U460 ( .A0(n114), .A1(n112), .B0(n113), .Y(n111) );
  OAI21XL U461 ( .A0(n114), .A1(n76), .B0(n77), .Y(n75) );
  INVX2 U462 ( .A(n81), .Y(n79) );
  OAI21X1 U463 ( .A0(n187), .A1(n185), .B0(n186), .Y(n184) );
  OAI21X1 U464 ( .A0(n199), .A1(n197), .B0(n198), .Y(n196) );
  AOI21X1 U465 ( .A0(n188), .A1(n196), .B0(n189), .Y(n187) );
  OAI21X1 U466 ( .A0(n190), .A1(n194), .B0(n191), .Y(n189) );
  NOR2X1 U467 ( .A(n193), .B(n190), .Y(n188) );
  OAI21XL U468 ( .A0(n133), .A1(n125), .B0(n128), .Y(n124) );
  NOR2X1 U469 ( .A(n132), .B(n125), .Y(n123) );
  CLKINVXL U470 ( .A(n131), .Y(n133) );
  XOR2X1 U471 ( .A(n122), .B(n11), .Y(SUM[29]) );
  XOR2X1 U472 ( .A(n129), .B(n12), .Y(SUM[28]) );
  NAND2X1 U473 ( .A(n268), .B(n128), .Y(n12) );
  INVX2 U474 ( .A(n211), .Y(n209) );
  AOI21X1 U475 ( .A0(n220), .A1(n431), .B0(n217), .Y(n215) );
  INVX2 U476 ( .A(n219), .Y(n217) );
  AOI21X1 U477 ( .A0(n204), .A1(n432), .B0(n201), .Y(n199) );
  INVX2 U478 ( .A(n203), .Y(n201) );
  AOI21X1 U479 ( .A0(n426), .A1(n240), .B0(n237), .Y(n235) );
  OAI21X1 U480 ( .A0(n205), .A1(n207), .B0(n206), .Y(n204) );
  OAI21X1 U481 ( .A0(n229), .A1(n231), .B0(n230), .Y(n228) );
  OAI21X1 U482 ( .A0(n221), .A1(n223), .B0(n222), .Y(n220) );
  OAI21X1 U483 ( .A0(n213), .A1(n215), .B0(n214), .Y(n212) );
  AOI21X1 U484 ( .A0(n228), .A1(n430), .B0(n225), .Y(n223) );
  INVX2 U485 ( .A(n227), .Y(n225) );
  OAI21X1 U486 ( .A0(n233), .A1(n235), .B0(n234), .Y(n232) );
  NAND2X1 U487 ( .A(n273), .B(n428), .Y(n150) );
  INVX2 U488 ( .A(n142), .Y(n140) );
  NOR2X1 U489 ( .A(n91), .B(n98), .Y(n89) );
  OAI21X1 U490 ( .A0(n91), .A1(n99), .B0(n92), .Y(n90) );
  AOI21X1 U491 ( .A0(n433), .A1(n425), .B0(n245), .Y(n243) );
  INVX2 U492 ( .A(n247), .Y(n245) );
  OAI21X1 U493 ( .A0(n241), .A1(n243), .B0(n242), .Y(n240) );
  INVX2 U494 ( .A(n44), .Y(n258) );
  OAI2BB1X1 U495 ( .A0N(n434), .A1N(n254), .B0(n253), .Y(n425) );
  CLKINVXL U496 ( .A(n80), .Y(n78) );
  CLKINVXL U497 ( .A(n60), .Y(n260) );
  XNOR2X1 U498 ( .A(n149), .B(n15), .Y(SUM[25]) );
  NAND2BX1 U499 ( .AN(n73), .B(n74), .Y(n5) );
  CLKINVXL U500 ( .A(n125), .Y(n268) );
  CLKINVXL U501 ( .A(n120), .Y(n267) );
  NAND2BX1 U502 ( .AN(n136), .B(n137), .Y(n13) );
  INVX2 U503 ( .A(n256), .Y(n254) );
  NAND2BX1 U504 ( .AN(n109), .B(n110), .Y(n9) );
  NAND2XL U505 ( .A(n273), .B(n158), .Y(n17) );
  NAND2X1 U506 ( .A(n429), .B(n171), .Y(n19) );
  XOR2XL U507 ( .A(n20), .B(n175), .Y(SUM[20]) );
  NAND2BX1 U508 ( .AN(n165), .B(n166), .Y(n18) );
  OAI21XL U509 ( .A0(n183), .A1(n181), .B0(n182), .Y(n180) );
  CLKINVXL U510 ( .A(n181), .Y(n278) );
  XOR2X1 U511 ( .A(n183), .B(n22), .Y(SUM[18]) );
  NAND2X1 U512 ( .A(n278), .B(n182), .Y(n22) );
  CLKINVXL U513 ( .A(n178), .Y(n277) );
  NAND2BX1 U514 ( .AN(n185), .B(n186), .Y(n23) );
  XOR2X1 U515 ( .A(n25), .B(n195), .Y(SUM[15]) );
  NAND2X1 U516 ( .A(n281), .B(n194), .Y(n25) );
  NAND2BX1 U517 ( .AN(n190), .B(n191), .Y(n24) );
  XOR2XL U518 ( .A(n26), .B(n199), .Y(SUM[14]) );
  NAND2X1 U519 ( .A(n432), .B(n203), .Y(n27) );
  NAND2BX1 U520 ( .AN(n205), .B(n206), .Y(n28) );
  XNOR2XL U521 ( .A(n29), .B(n212), .Y(SUM[11]) );
  NAND2X1 U522 ( .A(n427), .B(n211), .Y(n29) );
  NAND2BX1 U523 ( .AN(n221), .B(n222), .Y(n32) );
  XNOR2XL U524 ( .A(n33), .B(n228), .Y(SUM[7]) );
  NAND2X1 U525 ( .A(n430), .B(n227), .Y(n33) );
  XOR2XL U526 ( .A(n34), .B(n231), .Y(SUM[6]) );
  NAND2BX1 U527 ( .AN(n233), .B(n234), .Y(n35) );
  INVX2 U528 ( .A(n241), .Y(n293) );
  XOR2X1 U529 ( .A(n37), .B(n243), .Y(SUM[3]) );
  NAND2X1 U530 ( .A(n293), .B(n242), .Y(n37) );
  XNOR2X1 U531 ( .A(n38), .B(n425), .Y(SUM[2]) );
  NAND2X1 U532 ( .A(n433), .B(n247), .Y(n38) );
  NAND2X1 U533 ( .A(n434), .B(n253), .Y(n39) );
  XNOR2X1 U534 ( .A(n43), .B(n1), .Y(SUM[39]) );
  NOR2X1 U535 ( .A(B[37]), .B(A[37]), .Y(n53) );
  XNOR2X1 U536 ( .A(n111), .B(n9), .Y(SUM[31]) );
  XNOR2X1 U537 ( .A(n75), .B(n5), .Y(SUM[35]) );
  NOR2X1 U538 ( .A(B[25]), .B(A[25]), .Y(n147) );
  NOR2X1 U539 ( .A(B[14]), .B(A[14]), .Y(n197) );
  NOR2X1 U540 ( .A(B[20]), .B(A[20]), .Y(n173) );
  NOR2X1 U541 ( .A(B[26]), .B(A[26]), .Y(n141) );
  NOR2X1 U542 ( .A(B[16]), .B(A[16]), .Y(n190) );
  NOR2X1 U543 ( .A(B[31]), .B(A[31]), .Y(n109) );
  NAND2XL U544 ( .A(B[35]), .B(A[35]), .Y(n74) );
  NAND2XL U545 ( .A(B[36]), .B(A[36]), .Y(n63) );
  NOR2X1 U546 ( .A(B[23]), .B(A[23]), .Y(n157) );
  XOR2X1 U547 ( .A(n114), .B(n10), .Y(SUM[30]) );
  NOR2X1 U548 ( .A(B[10]), .B(A[10]), .Y(n213) );
  NOR2X1 U549 ( .A(B[15]), .B(A[15]), .Y(n193) );
  NAND2X1 U550 ( .A(B[26]), .B(A[26]), .Y(n142) );
  XOR2X1 U551 ( .A(n138), .B(n13), .Y(SUM[27]) );
  NOR2X1 U552 ( .A(B[12]), .B(A[12]), .Y(n205) );
  NOR2X1 U553 ( .A(B[17]), .B(A[17]), .Y(n185) );
  NOR2X1 U554 ( .A(B[5]), .B(A[5]), .Y(n233) );
  NOR2X1 U555 ( .A(B[32]), .B(A[32]), .Y(n98) );
  NOR2X1 U556 ( .A(B[6]), .B(A[6]), .Y(n229) );
  NAND2XL U557 ( .A(B[37]), .B(A[37]), .Y(n54) );
  NAND2XL U558 ( .A(B[27]), .B(A[27]), .Y(n137) );
  OR2XL U559 ( .A(B[9]), .B(A[9]), .Y(n431) );
  NAND2XL U560 ( .A(B[20]), .B(A[20]), .Y(n174) );
  NAND2XL U561 ( .A(B[14]), .B(A[14]), .Y(n198) );
  NOR2X1 U562 ( .A(B[33]), .B(A[33]), .Y(n91) );
  NAND2XL U563 ( .A(B[19]), .B(A[19]), .Y(n179) );
  NOR2X1 U564 ( .A(B[38]), .B(A[38]), .Y(n44) );
  NAND2XL U565 ( .A(B[24]), .B(A[24]), .Y(n155) );
  NAND2XL U566 ( .A(B[4]), .B(A[4]), .Y(n239) );
  OR2X1 U567 ( .A(B[2]), .B(A[2]), .Y(n433) );
  NAND2XL U568 ( .A(B[9]), .B(A[9]), .Y(n219) );
  NAND2XL U569 ( .A(B[5]), .B(A[5]), .Y(n234) );
  NOR2X1 U570 ( .A(B[3]), .B(A[3]), .Y(n241) );
  NAND2XL U571 ( .A(B[16]), .B(A[16]), .Y(n191) );
  NAND2XL U572 ( .A(B[10]), .B(A[10]), .Y(n214) );
  NAND2XL U573 ( .A(B[12]), .B(A[12]), .Y(n206) );
  NAND2X1 U574 ( .A(B[30]), .B(A[30]), .Y(n113) );
  NAND2XL U575 ( .A(B[29]), .B(A[29]), .Y(n121) );
  NOR2X1 U576 ( .A(B[8]), .B(A[8]), .Y(n221) );
  OR2XL U577 ( .A(B[1]), .B(A[1]), .Y(n434) );
  NAND2X1 U578 ( .A(B[38]), .B(A[39]), .Y(n42) );
  NOR2X1 U579 ( .A(B[38]), .B(A[39]), .Y(n41) );
  NAND2XL U580 ( .A(B[25]), .B(A[25]), .Y(n148) );
  NAND2XL U581 ( .A(B[6]), .B(A[6]), .Y(n230) );
  NAND2X1 U582 ( .A(B[32]), .B(A[32]), .Y(n99) );
  NAND2X1 U583 ( .A(B[38]), .B(A[38]), .Y(n45) );
  NAND2XL U584 ( .A(B[2]), .B(A[2]), .Y(n247) );
  NAND2XL U585 ( .A(B[1]), .B(A[1]), .Y(n253) );
  NAND2XL U586 ( .A(B[31]), .B(A[31]), .Y(n110) );
  NAND2XL U587 ( .A(B[3]), .B(A[3]), .Y(n242) );
  XNOR2X1 U588 ( .A(n143), .B(n14), .Y(SUM[26]) );
  NAND2XL U589 ( .A(B[33]), .B(A[33]), .Y(n92) );
  NOR2X1 U590 ( .A(B[22]), .B(A[22]), .Y(n165) );
  XOR2X1 U591 ( .A(n163), .B(n17), .Y(SUM[23]) );
  NAND2X1 U592 ( .A(B[0]), .B(A[0]), .Y(n256) );
  XNOR2X1 U593 ( .A(n192), .B(n24), .Y(SUM[16]) );
  XNOR2XL U594 ( .A(n27), .B(n204), .Y(SUM[13]) );
  XNOR2XL U595 ( .A(n31), .B(n220), .Y(SUM[9]) );
  XOR2XL U596 ( .A(n35), .B(n235), .Y(SUM[5]) );
  XNOR2X1 U597 ( .A(n36), .B(n240), .Y(SUM[4]) );
  XNOR2X1 U598 ( .A(n39), .B(n254), .Y(SUM[1]) );
  NAND2BX1 U599 ( .AN(n255), .B(n256), .Y(n40) );
  NOR2X1 U600 ( .A(B[0]), .B(A[0]), .Y(n255) );
  INVX2 U601 ( .A(n40), .Y(SUM[0]) );
  XOR2X1 U602 ( .A(n30), .B(n215), .Y(SUM[10]) );
  NOR2X1 U603 ( .A(n150), .B(n147), .Y(n145) );
  XOR2XL U604 ( .A(n18), .B(n167), .Y(SUM[22]) );
  XOR2XL U605 ( .A(n32), .B(n223), .Y(SUM[8]) );
  XNOR2X1 U606 ( .A(n172), .B(n19), .Y(SUM[21]) );
  XOR2XL U607 ( .A(n28), .B(n207), .Y(SUM[12]) );
  XOR2X1 U608 ( .A(n187), .B(n23), .Y(SUM[17]) );
  NOR2X1 U609 ( .A(n49), .B(n83), .Y(n47) );
endmodule


module MMSA_DW01_inc_10_DW01_inc_24 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  XOR2X1 U1 ( .A(carry[8]), .B(A[8]), .Y(SUM[8]) );
  CLKINVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module MMSA_DW01_inc_9_DW01_inc_23 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  CLKINVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module MMSA_DW01_inc_8_DW01_inc_22 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  ADDHXL U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  ADDHXL U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  ADDHXL U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADDHXL U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHXL U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  XOR2X1 U1 ( .A(carry[15]), .B(A[15]), .Y(SUM[15]) );
  CLKINVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module MMSA_DW01_inc_7_DW01_inc_21 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
  CLKINVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module MMSA_DW01_inc_6_DW01_inc_20 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  XOR2X1 U1 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
  CLKINVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module MMSA_DW01_inc_5_DW01_inc_19 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
  CLKINVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module MMSA_DW01_inc_4_DW01_inc_18 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  XOR2X1 U1 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
  CLKINVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module MMSA_DW01_inc_3_DW01_inc_17 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
  CLKINVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module MMSA_DW01_inc_2_DW01_inc_16 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
  CLKINVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module MMSA_DW01_inc_1_DW01_inc_15 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  XOR2X1 U1 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
  CLKINVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module MMSA_DW01_inc_0_DW01_inc_14 ( A, SUM );
  input [6:0] A;
  output [6:0] SUM;

  wire   [6:2] carry;

  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(carry[6]), .B(A[6]), .Y(SUM[6]) );
  CLKINVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module PE ( clk, rst, x_in0, x_in1, x_in2, x_in3, x_in4, x_in5, x_in6, x_in7, 
        w_in0, w_in1, w_in2, w_in3, w_in4, w_in5, w_in6, w_in7, y_out );
  input [15:0] x_in0;
  input [15:0] x_in1;
  input [15:0] x_in2;
  input [15:0] x_in3;
  input [15:0] x_in4;
  input [15:0] x_in5;
  input [15:0] x_in6;
  input [15:0] x_in7;
  input [15:0] w_in0;
  input [15:0] w_in1;
  input [15:0] w_in2;
  input [15:0] w_in3;
  input [15:0] w_in4;
  input [15:0] w_in5;
  input [15:0] w_in6;
  input [15:0] w_in7;
  output [39:0] y_out;
  input clk, rst;
  wire   N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N9, N89, N88, N87,
         N86, N85, N84, N83, N82, N81, N80, N8, N79, N78, N77, N76, N75, N74,
         N73, N72, N71, N70, N7, N69, N68, N67, N66, N65, N64, N63, N62, N61,
         N60, N6, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N5, N49,
         N48, N47, N468, N467, N466, N465, N464, N463, N462, N461, N460, N46,
         N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N45, N449,
         N448, N447, N446, N445, N444, N443, N442, N441, N440, N44, N439, N438,
         N437, N436, N435, N434, N433, N432, N431, N430, N43, N429, N428, N427,
         N426, N425, N424, N423, N422, N421, N420, N42, N419, N418, N417, N416,
         N415, N414, N413, N412, N411, N410, N41, N409, N408, N407, N406, N405,
         N404, N403, N402, N401, N400, N40, N4, N399, N398, N397, N396, N395,
         N394, N393, N392, N391, N390, N39, N389, N388, N387, N386, N385, N384,
         N383, N382, N381, N380, N38, N379, N378, N377, N376, N375, N374, N373,
         N372, N371, N370, N37, N369, N368, N367, N366, N365, N364, N363, N362,
         N361, N360, N36, N359, N358, N357, N356, N355, N354, N353, N352, N351,
         N350, N35, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340,
         N34, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N33,
         N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N32, N319,
         N318, N317, N316, N315, N314, N313, N312, N311, N310, N31, N309, N308,
         N307, N306, N305, N304, N303, N302, N301, N300, N30, N3, N299, N298,
         N297, N296, N295, N294, N293, N292, N291, N290, N29, N289, N288, N287,
         N286, N285, N284, N283, N282, N281, N280, N28, N279, N278, N277, N276,
         N275, N274, N273, N272, N271, N270, N27, N269, N268, N267, N266, N265,
         N264, N263, N262, N261, N260, N26, N259, N258, N257, N256, N255, N254,
         N253, N252, N251, N250, N25, N249, N248, N247, N246, N245, N244, N243,
         N242, N241, N240, N24, N239, N238, N237, N236, N235, N234, N233, N232,
         N231, N230, N23, N229, N228, N227, N226, N225, N224, N223, N222, N221,
         N220, N22, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210,
         N21, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N20,
         N2, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N19,
         N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N18, N179,
         N178, N177, N176, N175, N174, N173, N172, N171, N170, N17, N169, N168,
         N167, N166, N165, N164, N163, N162, N161, N160, N16, N159, N158, N157,
         N156, N155, N154, N153, N152, N151, N150, N15, N149, N148, N147, N146,
         N145, N144, N143, N142, N141, N140, N14, N139, N138, N137, N136, N135,
         N134, N133, N132, N131, N130, N13, N129, N128, N127, N126, N125, N124,
         N123, N122, N121, N120, N12, N119, N118, N117, N116, N115, N114, N113,
         N112, N111, N110, N11, N109, N108, N107, N106, N105, N104, N103, N102,
         N101, N100, N10, N1, N0, n1;

  PE_DW_mult_tc_19 mult_3077_6 ( .a(w_in5), .b(x_in5), .product({N329, N328, 
        N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, 
        N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, 
        N303, N302, N301, N300, N299, N298}) );
  PE_DW_mult_tc_16 mult_3077_8 ( .a(w_in7), .b(x_in7), .product({N468, N467, 
        N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, 
        N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, 
        N442, N441, N440, N439, N438, N437}) );
  PE_DW_mult_tc_22 mult_3077_5 ( .a(w_in4), .b(x_in4), .product({N261, N260, 
        N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, 
        N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, 
        N235, N234, N233, N232, N231, N230}) );
  PE_DW_mult_tc_17 mult_3077_7 ( .a(w_in6), .b(x_in6), .product({N398, N397, 
        N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, 
        N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, 
        N372, N371, N370, N369, N368, N367}) );
  PE_DW01_add_20 add_6_root_add_3077_7 ( .A({N31, N31, N30, N29, N28, N27, N26, 
        N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, 
        N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1, N0}), .B({N63, N63, N62, 
        N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, 
        N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, 
        N33, N32}), .CI(1'b0), .SUM({N96, N95, N94, N93, N92, N91, N90, N89, 
        N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, 
        N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64}) );
  PE_DW01_add_17 add_5_root_add_3077_7 ( .A({N128, N128, N128, N127, N126, 
        N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, 
        N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, 
        N101, N100, N99, N98, N97}), .B({N194, N194, N194, N193, N192, N191, 
        N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, 
        N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, 
        N166, N165, N164, N163}), .CI(1'b0), .SUM({N162, N161, N160, N159, 
        N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, 
        N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, 
        N134, N133, N132, N131, N130, N129}) );
  PE_DW01_add_23 add_0_root_add_3077_7 ( .A({N366, N366, N366, N365, N364, 
        N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, 
        N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, 
        N339, N338, N337, N336, N335, N334, N333, N332, N331, N330}), .B({N436, 
        N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, 
        N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, 
        N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, 
        N400, N399}), .CI(1'b0), .SUM(y_out[38:0]) );
  PE_DW01_add_22 add_1_root_add_3077_7 ( .A({N229, N229, N229, N229, N228, 
        N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, 
        N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, 
        N203, N202, N201, N200, N199, N198, N197, N196, N195}), .B({N297, N297, 
        N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, 
        N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, 
        N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262}), .CI(1'b0), .SUM({N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, 
        N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, 
        N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, 
        N402, N401, N400, N399}) );
  PE_DW01_add_21 add_4_root_add_3077_7 ( .A({N261, N261, N261, N261, N260, 
        N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, 
        N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, 
        N235, N234, N233, N232, N231, N230}), .B({N329, N329, N329, N329, N328, 
        N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, 
        N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, 
        N303, N302, N301, N300, N299, N298}), .CI(1'b0), .SUM({N229, N228, 
        N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, 
        N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, 
        N203, N202, N201, N200, N199, N198, N197, N196, N195}) );
  PE_DW01_add_24 add_3_root_add_3077_7 ( .A({N398, N398, N398, N398, N398, 
        N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, 
        N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, 
        N373, N372, N371, N370, N369, N368, N367}), .B({N468, N468, N468, N468, 
        N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, 
        N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, 
        N444, N443, N442, N441, N440, N439, N438, N437}), .CI(1'b0), .SUM({
        N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, 
        N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, 
        N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262}) );
  PE_DW01_add_26 add_2_root_add_3077_7 ( .A({N96, N96, N96, N96, N96, N95, N94, 
        N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, 
        N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, 
        N65, N64}), .B({N162, N162, N162, N162, N161, N160, N159, N158, N157, 
        N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, 
        N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, 
        N132, N131, N130, N129}), .CI(1'b0), .SUM({N366, N365, N364, N363, 
        N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, 
        N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, 
        N338, N337, N336, N335, N334, N333, N332, N331, N330}) );
  PE_DW_mult_tc_29 mult_3077_2 ( .a(w_in1), .b(x_in1), .product({N63, N62, N61, 
        N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, 
        N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, 
        N32}) );
  PE_DW_mult_tc_28 mult_3077 ( .a(w_in0), .b(x_in0), .product({N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2, N1, N0}) );
  PE_DW_mult_tc_31 mult_3077_4 ( .a(w_in3), .b(x_in3), .product({N194, N193, 
        N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, 
        N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, 
        N168, N167, N166, N165, N164, N163}) );
  PE_DW_mult_tc_30 mult_3077_3 ( .a(w_in2), .b(x_in2), .product({N128, N127, 
        N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, 
        N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, 
        N102, N101, N100, N99, N98, N97}) );
  INVX2 U1 ( .A(n1), .Y(y_out[39]) );
  CLKINVXL U2 ( .A(y_out[38]), .Y(n1) );
endmodule


module PE_DW_mult_tc_30 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n6, n9, n12, n16, n18, n22, n24, n28, n30, n34, n36, n40, n42, n46,
         n48, n51, n52, n53, n54, n55, n56, n58, n59, n60, n61, n63, n64, n66,
         n67, n68, n72, n73, n74, n75, n76, n77, n80, n82, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n103, n105, n106, n107, n108, n109, n110, n114, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n140, n141, n142,
         n143, n144, n145, n148, n149, n151, n154, n155, n156, n157, n158,
         n159, n160, n164, n166, n167, n168, n169, n170, n171, n173, n176,
         n177, n181, n182, n183, n184, n185, n186, n187, n188, n191, n192,
         n193, n194, n196, n199, n200, n201, n203, n204, n205, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n219, n220, n221,
         n222, n224, n227, n228, n229, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n244, n245, n246, n247, n248,
         n249, n251, n254, n255, n256, n257, n259, n261, n262, n264, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n281, n283, n284, n286, n288, n289, n290, n292, n294,
         n295, n296, n297, n298, n300, n302, n303, n304, n305, n307, n308,
         n311, n312, n313, n315, n316, n317, n319, n320, n323, n324, n325,
         n326, n329, n330, n336, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n844,
         n845, n846, n847, n848, n849, n850, n851, n867, n868, n869, n870,
         n871, n872, n874, n875, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980;

  AOI21X1 U56 ( .A0(n51), .A1(n85), .B0(n86), .Y(product[31]) );
  AOI21X1 U60 ( .A0(n123), .A1(n89), .B0(n90), .Y(n88) );
  AOI21X1 U68 ( .A0(n51), .A1(n94), .B0(n95), .Y(n93) );
  AOI21X1 U72 ( .A0(n123), .A1(n98), .B0(n99), .Y(n97) );
  AOI21X1 U76 ( .A0(n114), .A1(n970), .B0(n103), .Y(n101) );
  AOI21X1 U84 ( .A0(n51), .A1(n107), .B0(n108), .Y(n106) );
  AOI21X1 U88 ( .A0(n123), .A1(n969), .B0(n114), .Y(n110) );
  AOI21X1 U106 ( .A0(n126), .A1(n151), .B0(n127), .Y(n125) );
  AOI21X1 U114 ( .A0(n51), .A1(n131), .B0(n132), .Y(n130) );
  AOI21X1 U128 ( .A0(n51), .A1(n142), .B0(n143), .Y(n141) );
  AOI21X1 U132 ( .A0(n160), .A1(n313), .B0(n151), .Y(n145) );
  AOI21X1 U144 ( .A0(n51), .A1(n155), .B0(n156), .Y(n154) );
  AOI21X1 U160 ( .A0(n51), .A1(n168), .B0(n169), .Y(n167) );
  NAND2X4 U170 ( .A(n370), .B(n363), .Y(n171) );
  AOI21X1 U172 ( .A0(n51), .A1(n177), .B0(n960), .Y(n176) );
  NOR2X2 U181 ( .A(n378), .B(n371), .Y(n183) );
  AOI21X1 U184 ( .A0(n51), .A1(n186), .B0(n187), .Y(n185) );
  NOR2X2 U191 ( .A(n388), .B(n379), .Y(n188) );
  AOI21X1 U194 ( .A0(n51), .A1(n193), .B0(n194), .Y(n192) );
  OAI21X4 U214 ( .A0(n207), .A1(n235), .B0(n208), .Y(n51) );
  NOR2X2 U221 ( .A(n411), .B(n422), .Y(n211) );
  AOI21X1 U234 ( .A0(n234), .A1(n221), .B0(n222), .Y(n220) );
  OAI21X4 U240 ( .A0(n227), .A1(n233), .B0(n228), .Y(n222) );
  AOI21X1 U246 ( .A0(n234), .A1(n323), .B0(n231), .Y(n229) );
  NOR2X2 U251 ( .A(n451), .B(n464), .Y(n232) );
  NAND2X4 U252 ( .A(n451), .B(n464), .Y(n233) );
  NOR2X2 U256 ( .A(n241), .B(n238), .Y(n236) );
  OAI21X4 U284 ( .A0(n268), .A1(n256), .B0(n257), .Y(n255) );
  NOR2X2 U348 ( .A(n545), .B(n546), .Y(n296) );
  ADDFHX4 U381 ( .A(n367), .B(n365), .CI(n372), .CO(n362), .S(n363) );
  ADDFHX4 U385 ( .A(n382), .B(n373), .CI(n380), .CO(n370), .S(n371) );
  ADDFHX4 U388 ( .A(n972), .B(n580), .CI(n625), .CO(n376), .S(n377) );
  ADDFHX4 U394 ( .A(n402), .B(n400), .CI(n391), .CO(n388), .S(n389) );
  ADDFHX4 U401 ( .A(n420), .B(n405), .CI(n407), .CO(n402), .S(n403) );
  ADDFHX4 U405 ( .A(n415), .B(n424), .CI(n413), .CO(n410), .S(n411) );
  ADDFHX4 U408 ( .A(n629), .B(n614), .CI(n432), .CO(n416), .S(n417) );
  ADDFHX4 U411 ( .A(n427), .B(n438), .CI(n425), .CO(n422), .S(n423) );
  ADDFHX4 U418 ( .A(n441), .B(n452), .CI(n439), .CO(n436), .S(n437) );
  ADDFHX4 U419 ( .A(n456), .B(n443), .CI(n454), .CO(n438), .S(n439) );
  ADDFHX4 U426 ( .A(n455), .B(n466), .CI(n453), .CO(n450), .S(n451) );
  ADDFHX4 U427 ( .A(n461), .B(n457), .CI(n468), .CO(n452), .S(n453) );
  ADDFHX4 U439 ( .A(n481), .B(n490), .CI(n479), .CO(n476), .S(n477) );
  ADDFHX4 U445 ( .A(n493), .B(n500), .CI(n491), .CO(n488), .S(n489) );
  ADDFHX4 U446 ( .A(n504), .B(n502), .CI(n495), .CO(n490), .S(n491) );
  ADDFHX4 U450 ( .A(n503), .B(n510), .CI(n501), .CO(n498), .S(n499) );
  OAI22X1 U478 ( .A0(n48), .A1(n693), .B0(n46), .B1(n692), .Y(n338) );
  OAI22X1 U479 ( .A0(n48), .A1(n694), .B0(n46), .B1(n693), .Y(n565) );
  OAI22X1 U480 ( .A0(n48), .A1(n695), .B0(n46), .B1(n694), .Y(n344) );
  OAI22X1 U481 ( .A0(n48), .A1(n696), .B0(n46), .B1(n695), .Y(n566) );
  OAI22X1 U482 ( .A0(n48), .A1(n697), .B0(n46), .B1(n696), .Y(n354) );
  OAI22X1 U483 ( .A0(n48), .A1(n698), .B0(n46), .B1(n697), .Y(n567) );
  OAI22X1 U484 ( .A0(n48), .A1(n699), .B0(n46), .B1(n698), .Y(n368) );
  OAI22X1 U485 ( .A0(n48), .A1(n700), .B0(n46), .B1(n699), .Y(n568) );
  OAI22X1 U487 ( .A0(n48), .A1(n702), .B0(n46), .B1(n701), .Y(n569) );
  OAI22X1 U489 ( .A0(n48), .A1(n704), .B0(n46), .B1(n703), .Y(n570) );
  OAI22X1 U511 ( .A0(n42), .A1(n869), .B0(n40), .B1(n725), .Y(n557) );
  OAI22X1 U514 ( .A0(n42), .A1(n710), .B0(n709), .B1(n40), .Y(n575) );
  OAI22X1 U515 ( .A0(n42), .A1(n711), .B0(n710), .B1(n40), .Y(n576) );
  OAI22X1 U517 ( .A0(n42), .A1(n713), .B0(n712), .B1(n40), .Y(n578) );
  OAI22X1 U519 ( .A0(n42), .A1(n715), .B0(n714), .B1(n40), .Y(n580) );
  OAI22X1 U520 ( .A0(n42), .A1(n716), .B0(n715), .B1(n40), .Y(n581) );
  OAI22X1 U522 ( .A0(n42), .A1(n718), .B0(n717), .B1(n40), .Y(n583) );
  OAI22X1 U525 ( .A0(n42), .A1(n721), .B0(n720), .B1(n40), .Y(n586) );
  OAI22X1 U526 ( .A0(n42), .A1(n722), .B0(n721), .B1(n40), .Y(n587) );
  OAI22X1 U527 ( .A0(n42), .A1(n723), .B0(n722), .B1(n40), .Y(n588) );
  OAI22X1 U547 ( .A0(n36), .A1(n870), .B0(n34), .B1(n742), .Y(n558) );
  OAI22X1 U550 ( .A0(n36), .A1(n727), .B0(n726), .B1(n34), .Y(n592) );
  OAI22X1 U551 ( .A0(n36), .A1(n728), .B0(n727), .B1(n34), .Y(n593) );
  OAI22X1 U552 ( .A0(n36), .A1(n729), .B0(n728), .B1(n34), .Y(n594) );
  OAI22X1 U553 ( .A0(n36), .A1(n730), .B0(n729), .B1(n34), .Y(n595) );
  OAI22X1 U554 ( .A0(n36), .A1(n731), .B0(n730), .B1(n34), .Y(n596) );
  OAI22X1 U555 ( .A0(n36), .A1(n732), .B0(n731), .B1(n34), .Y(n597) );
  OAI22X1 U557 ( .A0(n36), .A1(n734), .B0(n733), .B1(n34), .Y(n599) );
  OAI22X1 U558 ( .A0(n36), .A1(n735), .B0(n734), .B1(n34), .Y(n600) );
  OAI22X1 U559 ( .A0(n36), .A1(n736), .B0(n735), .B1(n34), .Y(n601) );
  OAI22X1 U560 ( .A0(n36), .A1(n737), .B0(n736), .B1(n34), .Y(n602) );
  OAI22X1 U561 ( .A0(n36), .A1(n738), .B0(n737), .B1(n34), .Y(n603) );
  OAI22X1 U562 ( .A0(n36), .A1(n739), .B0(n738), .B1(n34), .Y(n604) );
  OAI22X1 U563 ( .A0(n36), .A1(n740), .B0(n739), .B1(n34), .Y(n605) );
  OAI22X1 U583 ( .A0(n30), .A1(n871), .B0(n28), .B1(n759), .Y(n559) );
  OAI22X1 U586 ( .A0(n30), .A1(n744), .B0(n743), .B1(n28), .Y(n609) );
  OAI22X1 U587 ( .A0(n30), .A1(n745), .B0(n744), .B1(n28), .Y(n610) );
  OAI22X1 U588 ( .A0(n30), .A1(n746), .B0(n745), .B1(n28), .Y(n611) );
  OAI22X1 U589 ( .A0(n30), .A1(n747), .B0(n746), .B1(n28), .Y(n612) );
  OAI22X1 U590 ( .A0(n30), .A1(n748), .B0(n747), .B1(n28), .Y(n613) );
  OAI22X1 U591 ( .A0(n30), .A1(n749), .B0(n748), .B1(n28), .Y(n614) );
  OAI22X1 U592 ( .A0(n30), .A1(n750), .B0(n749), .B1(n28), .Y(n615) );
  OAI22X1 U593 ( .A0(n30), .A1(n751), .B0(n750), .B1(n28), .Y(n616) );
  OAI22X1 U597 ( .A0(n30), .A1(n755), .B0(n754), .B1(n28), .Y(n620) );
  OAI22X1 U598 ( .A0(n30), .A1(n756), .B0(n755), .B1(n28), .Y(n621) );
  OAI22X1 U599 ( .A0(n30), .A1(n757), .B0(n756), .B1(n28), .Y(n622) );
  OAI22X1 U627 ( .A0(n24), .A1(n766), .B0(n765), .B1(n22), .Y(n631) );
  OAI22X1 U655 ( .A0(n18), .A1(n945), .B0(n16), .B1(n793), .Y(n561) );
  OAI22X1 U658 ( .A0(n18), .A1(n778), .B0(n777), .B1(n16), .Y(n643) );
  OAI22X1 U659 ( .A0(n18), .A1(n779), .B0(n778), .B1(n16), .Y(n644) );
  OAI22X1 U660 ( .A0(n18), .A1(n780), .B0(n779), .B1(n16), .Y(n645) );
  OAI22X1 U661 ( .A0(n18), .A1(n781), .B0(n780), .B1(n16), .Y(n646) );
  OAI22X1 U662 ( .A0(n18), .A1(n782), .B0(n781), .B1(n16), .Y(n647) );
  OAI22X1 U663 ( .A0(n18), .A1(n783), .B0(n782), .B1(n16), .Y(n648) );
  OAI22X1 U665 ( .A0(n18), .A1(n785), .B0(n784), .B1(n16), .Y(n650) );
  OAI22X1 U668 ( .A0(n18), .A1(n788), .B0(n787), .B1(n16), .Y(n653) );
  OAI22X1 U671 ( .A0(n18), .A1(n791), .B0(n790), .B1(n16), .Y(n656) );
  OAI22X1 U696 ( .A0(n12), .A1(n797), .B0(n796), .B1(n9), .Y(n662) );
  OAI22X1 U697 ( .A0(n12), .A1(n798), .B0(n797), .B1(n9), .Y(n663) );
  OAI22X1 U700 ( .A0(n12), .A1(n801), .B0(n800), .B1(n9), .Y(n666) );
  OAI22X1 U701 ( .A0(n12), .A1(n802), .B0(n801), .B1(n9), .Y(n667) );
  OAI22X1 U702 ( .A0(n12), .A1(n803), .B0(n802), .B1(n9), .Y(n668) );
  OAI22X1 U703 ( .A0(n12), .A1(n804), .B0(n803), .B1(n9), .Y(n669) );
  OAI22X1 U704 ( .A0(n12), .A1(n805), .B0(n804), .B1(n9), .Y(n670) );
  OAI22X1 U705 ( .A0(n12), .A1(n806), .B0(n805), .B1(n9), .Y(n671) );
  OAI22X1 U706 ( .A0(n12), .A1(n807), .B0(n806), .B1(n9), .Y(n672) );
  OAI22X1 U707 ( .A0(n12), .A1(n808), .B0(n807), .B1(n9), .Y(n673) );
  OAI22X1 U708 ( .A0(n12), .A1(n809), .B0(n808), .B1(n9), .Y(n674) );
  OAI22X1 U731 ( .A0(n6), .A1(n813), .B0(n812), .B1(n867), .Y(n678) );
  OAI22X1 U732 ( .A0(n6), .A1(n814), .B0(n813), .B1(n867), .Y(n679) );
  OAI22X1 U734 ( .A0(n6), .A1(n816), .B0(n815), .B1(n867), .Y(n681) );
  OAI22X1 U736 ( .A0(n6), .A1(n818), .B0(n817), .B1(n867), .Y(n683) );
  OAI22X1 U738 ( .A0(n6), .A1(n820), .B0(n819), .B1(n867), .Y(n685) );
  OAI22X1 U740 ( .A0(n6), .A1(n822), .B0(n821), .B1(n867), .Y(n687) );
  OAI22X1 U741 ( .A0(n6), .A1(n823), .B0(n822), .B1(n867), .Y(n688) );
  OAI22X1 U742 ( .A0(n6), .A1(n824), .B0(n823), .B1(n867), .Y(n689) );
  OAI22X1 U743 ( .A0(n6), .A1(n825), .B0(n824), .B1(n867), .Y(n690) );
  NAND2X4 U786 ( .A(n46), .B(n844), .Y(n48) );
  XNOR2X4 U788 ( .A(n979), .B(a[14]), .Y(n46) );
  NAND2X4 U789 ( .A(n40), .B(n845), .Y(n42) );
  XNOR2X4 U791 ( .A(n978), .B(a[12]), .Y(n40) );
  NAND2X4 U792 ( .A(n34), .B(n846), .Y(n36) );
  XNOR2X4 U794 ( .A(n977), .B(a[10]), .Y(n34) );
  NAND2X4 U795 ( .A(n28), .B(n847), .Y(n30) );
  XNOR2X4 U797 ( .A(n976), .B(a[8]), .Y(n28) );
  NAND2X4 U798 ( .A(n22), .B(n848), .Y(n24) );
  NAND2X4 U801 ( .A(n16), .B(n849), .Y(n18) );
  XNOR2X4 U803 ( .A(n974), .B(a[4]), .Y(n16) );
  NAND2X4 U804 ( .A(n9), .B(n850), .Y(n12) );
  XNOR2X4 U806 ( .A(n973), .B(a[2]), .Y(n9) );
  NAND2X4 U807 ( .A(n851), .B(n867), .Y(n6) );
  ADDHXL U812 ( .A(n679), .B(n649), .CO(n486), .S(n487) );
  BUFX12 U813 ( .A(a[13]), .Y(n979) );
  XOR2X4 U814 ( .A(n980), .B(a[14]), .Y(n844) );
  ADDFHX1 U815 ( .A(n557), .B(n664), .CI(n634), .CO(n484), .S(n485) );
  ADDFHX1 U816 ( .A(n635), .B(n665), .CI(n620), .CO(n494), .S(n495) );
  BUFX8 U817 ( .A(a[15]), .Y(n980) );
  NOR2X2 U818 ( .A(n477), .B(n488), .Y(n245) );
  XOR2X1 U819 ( .A(n176), .B(n61), .Y(product[23]) );
  XOR2X1 U820 ( .A(n220), .B(n67), .Y(product[17]) );
  XOR2X1 U821 ( .A(n117), .B(n56), .Y(product[28]) );
  XOR2X1 U822 ( .A(n106), .B(n55), .Y(product[29]) );
  XOR2X1 U823 ( .A(n167), .B(n60), .Y(product[24]) );
  XOR2X1 U824 ( .A(n154), .B(n59), .Y(product[25]) );
  XOR2X1 U825 ( .A(n141), .B(n58), .Y(product[26]) );
  XNOR2X1 U826 ( .A(n130), .B(n956), .Y(product[27]) );
  XOR2X1 U827 ( .A(n201), .B(n64), .Y(product[20]) );
  ADDFX2 U828 ( .A(n569), .B(n582), .CI(n612), .CO(n394), .S(n395) );
  ADDFX2 U829 ( .A(n567), .B(n593), .CI(n366), .CO(n358), .S(n359) );
  ADDFHX1 U830 ( .A(n616), .B(n971), .CI(n676), .CO(n446), .S(n447) );
  NOR2X1 U831 ( .A(n356), .B(n351), .Y(n148) );
  CMPR32X1 U832 ( .A(n361), .B(n359), .C(n364), .CO(n356), .S(n357) );
  CLKINVXL U833 ( .A(n158), .Y(n160) );
  NOR2X1 U834 ( .A(n148), .B(n137), .Y(n135) );
  NAND2X1 U835 ( .A(n159), .B(n135), .Y(n133) );
  ADDFX2 U836 ( .A(n360), .B(n353), .CI(n358), .CO(n350), .S(n351) );
  ADDFX2 U837 ( .A(n566), .B(n352), .CI(n349), .CO(n346), .S(n347) );
  ADDFHX1 U838 ( .A(n392), .B(n390), .CI(n381), .CO(n378), .S(n379) );
  NAND2X2 U839 ( .A(n489), .B(n498), .Y(n249) );
  NAND2X1 U840 ( .A(n477), .B(n488), .Y(n246) );
  NOR2X1 U841 ( .A(n350), .B(n347), .Y(n137) );
  NAND2X1 U842 ( .A(n399), .B(n410), .Y(n205) );
  NAND2XL U843 ( .A(n411), .B(n422), .Y(n212) );
  OAI21X2 U844 ( .A0(n242), .A1(n238), .B0(n239), .Y(n237) );
  NOR2X2 U845 ( .A(n423), .B(n436), .Y(n216) );
  OAI21X1 U846 ( .A0(n211), .A1(n219), .B0(n212), .Y(n210) );
  NOR2X1 U847 ( .A(n6), .B(n819), .Y(n949) );
  NOR2X1 U848 ( .A(n818), .B(n867), .Y(n950) );
  OAI22X2 U849 ( .A0(n6), .A1(n821), .B0(n820), .B1(n867), .Y(n686) );
  XOR2X1 U850 ( .A(n80), .B(n298), .Y(product[4]) );
  ADDFX2 U851 ( .A(n596), .B(n626), .CI(n387), .CO(n384), .S(n385) );
  ADDFX2 U852 ( .A(n636), .B(n621), .CI(n507), .CO(n502), .S(n503) );
  ADDFX2 U853 ( .A(n618), .B(n663), .CI(n648), .CO(n472), .S(n473) );
  ADDFX2 U854 ( .A(n633), .B(n603), .CI(n486), .CO(n470), .S(n471) );
  ADDFX2 U855 ( .A(n619), .B(n589), .CI(n604), .CO(n482), .S(n483) );
  ADDFX2 U856 ( .A(n594), .B(n579), .CI(n369), .CO(n366), .S(n367) );
  ADDFX2 U857 ( .A(n609), .B(n376), .CI(n374), .CO(n364), .S(n365) );
  XOR2X1 U858 ( .A(n247), .B(n955), .Y(product[13]) );
  ADDFX2 U859 ( .A(n592), .B(n577), .CI(n355), .CO(n352), .S(n353) );
  ADDFX2 U860 ( .A(n611), .B(n581), .CI(n396), .CO(n382), .S(n383) );
  ADDFX2 U861 ( .A(n384), .B(n377), .CI(n375), .CO(n372), .S(n373) );
  ADDFX2 U862 ( .A(n394), .B(n385), .CI(n383), .CO(n380), .S(n381) );
  ADDFX2 U863 ( .A(n627), .B(n406), .CI(n404), .CO(n392), .S(n393) );
  ADDFHX1 U864 ( .A(n395), .B(n397), .CI(n393), .CO(n390), .S(n391) );
  ADDFX2 U865 ( .A(n418), .B(n416), .CI(n414), .CO(n400), .S(n401) );
  OAI21X1 U866 ( .A0(n278), .A1(n290), .B0(n279), .Y(n277) );
  AOI21X1 U867 ( .A0(n964), .A1(n286), .B0(n281), .Y(n279) );
  NOR2X1 U868 ( .A(n489), .B(n498), .Y(n248) );
  ADDFX2 U869 ( .A(n487), .B(n496), .CI(n494), .CO(n480), .S(n481) );
  ADDFX2 U870 ( .A(n434), .B(n599), .CI(n659), .CO(n420), .S(n421) );
  ADDFHX1 U871 ( .A(n662), .B(n463), .CI(n474), .CO(n456), .S(n457) );
  ADDFX2 U872 ( .A(n645), .B(n585), .CI(n630), .CO(n430), .S(n431) );
  OAI22X1 U873 ( .A0(n12), .A1(n795), .B0(n794), .B1(n9), .Y(n660) );
  ADDFHX1 U874 ( .A(n462), .B(n449), .CI(n460), .CO(n442), .S(n443) );
  XNOR2X1 U875 ( .A(n631), .B(n571), .Y(n449) );
  ADDFX2 U876 ( .A(n600), .B(n448), .CI(n446), .CO(n428), .S(n429) );
  ADDFX2 U877 ( .A(n475), .B(n484), .CI(n473), .CO(n468), .S(n469) );
  CMPR32X1 U878 ( .A(n472), .B(n470), .C(n459), .CO(n454), .S(n455) );
  ADDFX2 U879 ( .A(n482), .B(n471), .CI(n480), .CO(n466), .S(n467) );
  ADDFHX1 U880 ( .A(n403), .B(n412), .CI(n401), .CO(n398), .S(n399) );
  CMPR32X1 U881 ( .A(n430), .B(n421), .C(n419), .CO(n414), .S(n415) );
  ADDFX2 U882 ( .A(n458), .B(n447), .CI(n445), .CO(n440), .S(n441) );
  ADDFHX1 U883 ( .A(n442), .B(n429), .CI(n440), .CO(n424), .S(n425) );
  ADDFX2 U884 ( .A(n469), .B(n478), .CI(n467), .CO(n464), .S(n465) );
  INVX2 U885 ( .A(a[0]), .Y(n867) );
  NAND2X1 U886 ( .A(n122), .B(n969), .Y(n109) );
  NOR2X1 U887 ( .A(n370), .B(n363), .Y(n170) );
  OAI21X1 U888 ( .A0(n52), .A1(n133), .B0(n134), .Y(n132) );
  AOI21X1 U889 ( .A0(n160), .A1(n135), .B0(n136), .Y(n134) );
  NOR2X1 U890 ( .A(n53), .B(n133), .Y(n131) );
  NAND2X1 U891 ( .A(n320), .B(n212), .Y(n66) );
  NOR2X1 U892 ( .A(n346), .B(n343), .Y(n128) );
  NOR2X1 U893 ( .A(n137), .B(n128), .Y(n126) );
  AOI21X1 U894 ( .A0(n962), .A1(n173), .B0(n164), .Y(n158) );
  INVX2 U895 ( .A(n171), .Y(n173) );
  NOR2X1 U896 ( .A(n399), .B(n410), .Y(n204) );
  NOR2X2 U897 ( .A(n465), .B(n476), .Y(n238) );
  NAND2X1 U898 ( .A(n325), .B(n326), .Y(n241) );
  INVX2 U899 ( .A(n246), .Y(n244) );
  INVX2 U900 ( .A(n249), .Y(n251) );
  INVX2 U901 ( .A(n182), .Y(n961) );
  OAI21X1 U902 ( .A0(n183), .A1(n191), .B0(n184), .Y(n182) );
  NOR2X1 U903 ( .A(n188), .B(n183), .Y(n181) );
  NOR2X1 U904 ( .A(n204), .B(n199), .Y(n193) );
  NOR2X1 U905 ( .A(n157), .B(n124), .Y(n122) );
  NAND2X1 U906 ( .A(n193), .B(n181), .Y(n53) );
  NAND2X1 U907 ( .A(n209), .B(n221), .Y(n207) );
  OAI22X1 U908 ( .A0(n24), .A1(n772), .B0(n771), .B1(n22), .Y(n637) );
  NOR2BX1 U909 ( .AN(b[0]), .B(n22), .Y(n641) );
  OAI22XL U910 ( .A0(n24), .A1(n775), .B0(n774), .B1(n22), .Y(n640) );
  OAI22X1 U911 ( .A0(n24), .A1(n872), .B0(n22), .B1(n776), .Y(n560) );
  OAI22X1 U912 ( .A0(n12), .A1(n799), .B0(n798), .B1(n9), .Y(n664) );
  OAI22X2 U913 ( .A0(n6), .A1(n815), .B0(n814), .B1(n867), .Y(n680) );
  OR2X2 U914 ( .A(n499), .B(n508), .Y(n943) );
  OR2X1 U915 ( .A(n691), .B(n563), .Y(n944) );
  INVX2 U916 ( .A(n960), .Y(n52) );
  OAI2BB1X1 U917 ( .A0N(n194), .A1N(n181), .B0(n961), .Y(n960) );
  BUFX8 U918 ( .A(a[5]), .Y(n975) );
  INVX2 U919 ( .A(n975), .Y(n945) );
  AOI21X2 U920 ( .A0(n943), .A1(n264), .B0(n259), .Y(n257) );
  OAI21X1 U921 ( .A0(n254), .A1(n248), .B0(n249), .Y(n247) );
  OAI22X2 U922 ( .A0(n18), .A1(n787), .B0(n786), .B1(n16), .Y(n652) );
  AOI21XL U923 ( .A0(n214), .A1(n234), .B0(n215), .Y(n213) );
  ADDFHX1 U924 ( .A(n607), .B(n682), .CI(n622), .CO(n514), .S(n515) );
  OAI21X1 U925 ( .A0(n254), .A1(n241), .B0(n242), .Y(n240) );
  OAI22X2 U926 ( .A0(n6), .A1(n817), .B0(n816), .B1(n867), .Y(n682) );
  NAND2X2 U927 ( .A(n975), .B(a[6]), .Y(n947) );
  NAND2X4 U928 ( .A(n945), .B(n946), .Y(n948) );
  NAND2X4 U929 ( .A(n947), .B(n948), .Y(n22) );
  INVX2 U930 ( .A(a[6]), .Y(n946) );
  OAI22XL U931 ( .A0(n24), .A1(n774), .B0(n773), .B1(n22), .Y(n639) );
  OAI22XL U932 ( .A0(n24), .A1(n769), .B0(n768), .B1(n22), .Y(n634) );
  OAI22XL U933 ( .A0(n24), .A1(n768), .B0(n767), .B1(n22), .Y(n633) );
  OAI22XL U934 ( .A0(n24), .A1(n765), .B0(n764), .B1(n22), .Y(n630) );
  OAI22XL U935 ( .A0(n24), .A1(n763), .B0(n762), .B1(n22), .Y(n628) );
  OAI22XL U936 ( .A0(n24), .A1(n762), .B0(n761), .B1(n22), .Y(n627) );
  OAI22XL U937 ( .A0(n24), .A1(n770), .B0(n769), .B1(n22), .Y(n635) );
  OAI22XL U938 ( .A0(n24), .A1(n771), .B0(n770), .B1(n22), .Y(n636) );
  OAI22XL U939 ( .A0(n24), .A1(n773), .B0(n772), .B1(n22), .Y(n638) );
  OAI22XL U940 ( .A0(n24), .A1(n767), .B0(n766), .B1(n22), .Y(n632) );
  OAI22XL U941 ( .A0(n24), .A1(n764), .B0(n763), .B1(n22), .Y(n629) );
  OR2X2 U942 ( .A(n949), .B(n950), .Y(n684) );
  ADDFHX1 U943 ( .A(n624), .B(n684), .CI(n639), .CO(n528), .S(n529) );
  INVXL U944 ( .A(n235), .Y(n234) );
  AOI21X2 U945 ( .A0(n269), .A1(n277), .B0(n270), .Y(n268) );
  CMPR32X1 U946 ( .A(n521), .B(n526), .C(n519), .CO(n516), .S(n517) );
  INVX3 U947 ( .A(n255), .Y(n254) );
  NOR2X1 U948 ( .A(n227), .B(n232), .Y(n221) );
  OR2X2 U949 ( .A(n509), .B(n516), .Y(n963) );
  NOR2X1 U950 ( .A(n525), .B(n530), .Y(n274) );
  XOR2X1 U951 ( .A(n959), .B(n303), .Y(product[3]) );
  AND2X1 U952 ( .A(n316), .B(n184), .Y(n954) );
  NAND2X1 U953 ( .A(n509), .B(n516), .Y(n266) );
  ADDFX1 U954 ( .A(n561), .B(n672), .CI(n543), .CO(n540), .S(n541) );
  XOR2X1 U955 ( .A(n973), .B(a[0]), .Y(n851) );
  XNOR2X1 U956 ( .A(n980), .B(b[8]), .Y(n699) );
  AOI21XL U957 ( .A0(n51), .A1(n319), .B0(n203), .Y(n201) );
  NAND2X1 U958 ( .A(n465), .B(n476), .Y(n239) );
  XNOR2X1 U959 ( .A(n185), .B(n954), .Y(product[22]) );
  CLKINVXL U960 ( .A(n148), .Y(n313) );
  AND2X1 U961 ( .A(n311), .B(n129), .Y(n956) );
  NAND2XL U962 ( .A(n378), .B(n371), .Y(n184) );
  NAND2X1 U963 ( .A(n388), .B(n379), .Y(n191) );
  OR2X4 U964 ( .A(n531), .B(n536), .Y(n964) );
  ADDFHX1 U965 ( .A(n559), .B(n623), .CI(n638), .CO(n520), .S(n521) );
  NAND2BXL U966 ( .AN(b[0]), .B(n976), .Y(n776) );
  CLKINVXL U967 ( .A(n354), .Y(n355) );
  BUFX20 U968 ( .A(a[1]), .Y(n973) );
  BUFX20 U969 ( .A(a[7]), .Y(n976) );
  BUFX20 U970 ( .A(a[3]), .Y(n974) );
  BUFX20 U971 ( .A(a[9]), .Y(n977) );
  BUFX20 U972 ( .A(a[11]), .Y(n978) );
  OAI21X2 U973 ( .A0(n199), .A1(n205), .B0(n200), .Y(n194) );
  XOR2X1 U974 ( .A(n240), .B(n951), .Y(product[14]) );
  AND2X2 U975 ( .A(n324), .B(n239), .Y(n951) );
  NAND2BX1 U976 ( .AN(n199), .B(n200), .Y(n64) );
  OAI21XL U977 ( .A0(n52), .A1(n157), .B0(n158), .Y(n156) );
  XOR2X1 U978 ( .A(n234), .B(n952), .Y(product[15]) );
  AND2X1 U979 ( .A(n323), .B(n233), .Y(n952) );
  XOR2X1 U980 ( .A(n51), .B(n953), .Y(product[19]) );
  AND2X1 U981 ( .A(n319), .B(n205), .Y(n953) );
  OAI21XL U982 ( .A0(n52), .A1(n144), .B0(n145), .Y(n143) );
  NAND2BX1 U983 ( .AN(n216), .B(n219), .Y(n67) );
  NAND2BX1 U984 ( .AN(n227), .B(n228), .Y(n68) );
  XOR2X1 U985 ( .A(n213), .B(n66), .Y(product[18]) );
  NAND2XL U986 ( .A(n159), .B(n313), .Y(n144) );
  NAND2X1 U987 ( .A(n389), .B(n398), .Y(n200) );
  NAND2XL U988 ( .A(n962), .B(n166), .Y(n60) );
  AND2X1 U989 ( .A(n325), .B(n246), .Y(n955) );
  CLKINVXL U990 ( .A(n53), .Y(n177) );
  INVX2 U991 ( .A(n248), .Y(n326) );
  NAND2X1 U992 ( .A(n423), .B(n436), .Y(n219) );
  CLKINVXL U993 ( .A(n188), .Y(n317) );
  NAND2XL U994 ( .A(n313), .B(n149), .Y(n59) );
  XNOR2X1 U995 ( .A(n267), .B(n74), .Y(product[10]) );
  XOR2X1 U996 ( .A(n262), .B(n73), .Y(product[11]) );
  AOI21XL U997 ( .A0(n267), .A1(n963), .B0(n264), .Y(n262) );
  INVX2 U998 ( .A(n170), .Y(n315) );
  XOR2X1 U999 ( .A(n276), .B(n76), .Y(product[8]) );
  CLKINVXL U1000 ( .A(n277), .Y(n276) );
  XNOR2X1 U1001 ( .A(n273), .B(n75), .Y(product[9]) );
  NAND2XL U1002 ( .A(n329), .B(n272), .Y(n75) );
  CLKINVXL U1003 ( .A(n271), .Y(n329) );
  NAND2X1 U1004 ( .A(n313), .B(n126), .Y(n124) );
  OAI21X1 U1005 ( .A0(n149), .A1(n137), .B0(n140), .Y(n136) );
  NAND2XL U1006 ( .A(n499), .B(n508), .Y(n261) );
  AOI21X1 U1007 ( .A0(n295), .A1(n966), .B0(n292), .Y(n290) );
  CLKINVX2 U1008 ( .A(n294), .Y(n292) );
  NAND2XL U1009 ( .A(n525), .B(n530), .Y(n275) );
  INVX1 U1010 ( .A(n288), .Y(n286) );
  NAND2XL U1011 ( .A(n312), .B(n140), .Y(n58) );
  XOR2X1 U1012 ( .A(n957), .B(n289), .Y(product[6]) );
  AND2X1 U1013 ( .A(n967), .B(n288), .Y(n957) );
  NAND2XL U1014 ( .A(n362), .B(n357), .Y(n166) );
  XNOR2XL U1015 ( .A(n958), .B(n295), .Y(product[5]) );
  NAND2XL U1016 ( .A(n966), .B(n294), .Y(n958) );
  XOR2X1 U1017 ( .A(n284), .B(n77), .Y(product[7]) );
  AOI21XL U1018 ( .A0(n289), .A1(n967), .B0(n286), .Y(n284) );
  NAND2BX1 U1019 ( .AN(n296), .B(n297), .Y(n80) );
  AND2X1 U1020 ( .A(n965), .B(n302), .Y(n959) );
  XOR2XL U1021 ( .A(n82), .B(n307), .Y(product[2]) );
  NAND2XL U1022 ( .A(n336), .B(n305), .Y(n82) );
  CLKINVXL U1023 ( .A(n304), .Y(n336) );
  OAI21XL U1024 ( .A0(n140), .A1(n128), .B0(n129), .Y(n127) );
  OAI21XL U1025 ( .A0(n158), .A1(n124), .B0(n125), .Y(n123) );
  ADDFHX2 U1026 ( .A(n428), .B(n417), .CI(n426), .CO(n412), .S(n413) );
  ADDFHX1 U1027 ( .A(n522), .B(n515), .CI(n520), .CO(n510), .S(n511) );
  NAND2XL U1028 ( .A(n531), .B(n536), .Y(n283) );
  NAND2XL U1029 ( .A(n547), .B(n674), .Y(n302) );
  INVX2 U1030 ( .A(n434), .Y(n435) );
  ADDFHX1 U1031 ( .A(n615), .B(n660), .CI(n435), .CO(n432), .S(n433) );
  ADDFHX1 U1032 ( .A(n590), .B(n680), .CI(n605), .CO(n496), .S(n497) );
  CLKINVXL U1033 ( .A(n794), .Y(n554) );
  ADDFX1 U1034 ( .A(n573), .B(n678), .CI(n588), .CO(n474), .S(n475) );
  OAI22XL U1035 ( .A0(n42), .A1(n720), .B0(n719), .B1(n40), .Y(n585) );
  OAI22XL U1036 ( .A0(n42), .A1(n717), .B0(n716), .B1(n40), .Y(n582) );
  OAI22XL U1037 ( .A0(n36), .A1(n733), .B0(n732), .B1(n34), .Y(n598) );
  OAI22XL U1038 ( .A0(n18), .A1(n789), .B0(n788), .B1(n16), .Y(n654) );
  OAI22XL U1039 ( .A0(n30), .A1(n754), .B0(n753), .B1(n28), .Y(n619) );
  ADDFX1 U1040 ( .A(n671), .B(n542), .CI(n539), .CO(n536), .S(n537) );
  OAI22XL U1041 ( .A0(n12), .A1(n874), .B0(n9), .B1(n810), .Y(n562) );
  OAI22XL U1042 ( .A0(n18), .A1(n790), .B0(n789), .B1(n16), .Y(n655) );
  ADDHXL U1043 ( .A(n677), .B(n647), .CO(n462), .S(n463) );
  OAI22XL U1044 ( .A0(n6), .A1(n812), .B0(n811), .B1(n867), .Y(n677) );
  OAI22XL U1045 ( .A0(n12), .A1(n800), .B0(n799), .B1(n9), .Y(n665) );
  ADDHXL U1046 ( .A(n681), .B(n651), .CO(n506), .S(n507) );
  OAI22XL U1047 ( .A0(n18), .A1(n786), .B0(n785), .B1(n16), .Y(n651) );
  OAI22XL U1048 ( .A0(n24), .A1(n761), .B0(n760), .B1(n22), .Y(n626) );
  XNOR2X1 U1049 ( .A(b[0]), .B(n980), .Y(n707) );
  OAI22XL U1050 ( .A0(n36), .A1(n741), .B0(n740), .B1(n34), .Y(n606) );
  OAI22XL U1051 ( .A0(n42), .A1(n719), .B0(n718), .B1(n40), .Y(n584) );
  OAI22XL U1052 ( .A0(n18), .A1(n784), .B0(n783), .B1(n16), .Y(n649) );
  OAI22XL U1053 ( .A0(n42), .A1(n714), .B0(n713), .B1(n40), .Y(n579) );
  NAND2BX1 U1054 ( .AN(b[0]), .B(n978), .Y(n742) );
  OAI22XL U1055 ( .A0(n42), .A1(n712), .B0(n711), .B1(n40), .Y(n577) );
  CLKINVXL U1056 ( .A(n811), .Y(n555) );
  CLKINVXL U1057 ( .A(n726), .Y(n550) );
  ADDFX1 U1058 ( .A(n354), .B(n576), .CI(n591), .CO(n348), .S(n349) );
  XOR2X1 U1059 ( .A(n977), .B(a[8]), .Y(n847) );
  XNOR2X1 U1060 ( .A(n980), .B(b[3]), .Y(n704) );
  XNOR2X1 U1061 ( .A(n980), .B(b[2]), .Y(n705) );
  XNOR2X1 U1062 ( .A(n975), .B(b[15]), .Y(n777) );
  XNOR2X1 U1063 ( .A(n980), .B(b[4]), .Y(n703) );
  XNOR2X1 U1064 ( .A(n980), .B(b[6]), .Y(n701) );
  XNOR2X1 U1065 ( .A(n980), .B(b[7]), .Y(n700) );
  XNOR2X1 U1066 ( .A(n980), .B(b[9]), .Y(n698) );
  XNOR2X1 U1067 ( .A(n980), .B(b[10]), .Y(n697) );
  XNOR2X1 U1068 ( .A(n977), .B(b[15]), .Y(n743) );
  XNOR2X1 U1069 ( .A(n980), .B(b[11]), .Y(n696) );
  XNOR2X1 U1070 ( .A(n980), .B(b[12]), .Y(n695) );
  XNOR2X1 U1071 ( .A(n980), .B(b[13]), .Y(n694) );
  XNOR2X1 U1072 ( .A(n980), .B(b[14]), .Y(n693) );
  XNOR2X1 U1073 ( .A(n980), .B(b[15]), .Y(n692) );
  INVX2 U1074 ( .A(n122), .Y(n120) );
  NOR2X1 U1075 ( .A(n53), .B(n144), .Y(n142) );
  NOR2X1 U1076 ( .A(n53), .B(n96), .Y(n94) );
  NOR2X2 U1077 ( .A(n211), .B(n216), .Y(n209) );
  CLKINVXL U1078 ( .A(n211), .Y(n320) );
  NOR2BXL U1079 ( .AN(n221), .B(n216), .Y(n214) );
  OAI21XL U1080 ( .A0(n224), .A1(n216), .B0(n219), .Y(n215) );
  CLKINVXL U1081 ( .A(n222), .Y(n224) );
  INVX2 U1082 ( .A(n268), .Y(n267) );
  INVX2 U1083 ( .A(n157), .Y(n159) );
  CLKINVXL U1084 ( .A(n238), .Y(n324) );
  CLKINVXL U1085 ( .A(n204), .Y(n319) );
  CLKINVXL U1086 ( .A(n232), .Y(n323) );
  CLKINVXL U1087 ( .A(n205), .Y(n203) );
  CLKINVXL U1088 ( .A(n233), .Y(n231) );
  NAND2XL U1089 ( .A(n122), .B(n98), .Y(n96) );
  XOR2X2 U1090 ( .A(n192), .B(n63), .Y(product[21]) );
  NAND2X1 U1091 ( .A(n317), .B(n191), .Y(n63) );
  NAND2XL U1092 ( .A(n315), .B(n171), .Y(n61) );
  NOR2XL U1093 ( .A(n53), .B(n157), .Y(n155) );
  NAND2X2 U1094 ( .A(n437), .B(n450), .Y(n228) );
  NAND2X2 U1095 ( .A(n943), .B(n963), .Y(n256) );
  INVX2 U1096 ( .A(n261), .Y(n259) );
  OAI21X1 U1097 ( .A0(n271), .A1(n275), .B0(n272), .Y(n270) );
  NOR2X1 U1098 ( .A(n271), .B(n274), .Y(n269) );
  OAI21XL U1099 ( .A0(n52), .A1(n170), .B0(n171), .Y(n169) );
  NOR2XL U1100 ( .A(n53), .B(n170), .Y(n168) );
  OAI21XL U1101 ( .A0(n52), .A1(n120), .B0(n121), .Y(n119) );
  INVX2 U1102 ( .A(n123), .Y(n121) );
  NAND2X1 U1103 ( .A(n315), .B(n962), .Y(n157) );
  INVX2 U1104 ( .A(n166), .Y(n164) );
  CLKINVXL U1105 ( .A(n183), .Y(n316) );
  NAND2X1 U1106 ( .A(n963), .B(n266), .Y(n74) );
  INVX2 U1107 ( .A(n266), .Y(n264) );
  INVX2 U1108 ( .A(n290), .Y(n289) );
  NAND2X1 U1109 ( .A(n330), .B(n275), .Y(n76) );
  INVX2 U1110 ( .A(n274), .Y(n330) );
  XOR2X1 U1111 ( .A(n254), .B(n72), .Y(product[12]) );
  NAND2XL U1112 ( .A(n326), .B(n249), .Y(n72) );
  NOR2BXL U1113 ( .AN(n193), .B(n188), .Y(n186) );
  NAND2XL U1114 ( .A(n943), .B(n261), .Y(n73) );
  OAI21X1 U1115 ( .A0(n276), .A1(n274), .B0(n275), .Y(n273) );
  CLKINVXL U1116 ( .A(n194), .Y(n196) );
  INVX2 U1117 ( .A(n149), .Y(n151) );
  OAI21XL U1118 ( .A0(n52), .A1(n96), .B0(n97), .Y(n95) );
  INVX2 U1119 ( .A(n101), .Y(n99) );
  NAND2XL U1120 ( .A(n122), .B(n89), .Y(n87) );
  OAI21XL U1121 ( .A0(n52), .A1(n87), .B0(n88), .Y(n86) );
  NOR2X1 U1122 ( .A(n53), .B(n87), .Y(n85) );
  INVX2 U1123 ( .A(n100), .Y(n98) );
  INVX2 U1124 ( .A(n128), .Y(n311) );
  CLKINVXL U1125 ( .A(n137), .Y(n312) );
  NAND2X1 U1126 ( .A(n964), .B(n967), .Y(n278) );
  INVX2 U1127 ( .A(n283), .Y(n281) );
  NAND2X1 U1128 ( .A(n969), .B(n116), .Y(n56) );
  NOR2XL U1129 ( .A(n53), .B(n120), .Y(n118) );
  OAI21XL U1130 ( .A0(n52), .A1(n109), .B0(n110), .Y(n108) );
  NAND2X1 U1131 ( .A(n970), .B(n105), .Y(n55) );
  NOR2X1 U1132 ( .A(n517), .B(n524), .Y(n271) );
  OR2X4 U1133 ( .A(n362), .B(n357), .Y(n962) );
  AOI21X1 U1134 ( .A0(n965), .A1(n303), .B0(n300), .Y(n298) );
  INVX2 U1135 ( .A(n302), .Y(n300) );
  OAI21XL U1136 ( .A0(n298), .A1(n296), .B0(n297), .Y(n295) );
  NAND2X1 U1137 ( .A(n517), .B(n524), .Y(n272) );
  NAND2X1 U1138 ( .A(n964), .B(n283), .Y(n77) );
  NAND2X1 U1139 ( .A(n356), .B(n351), .Y(n149) );
  XOR2X1 U1140 ( .A(n93), .B(n54), .Y(product[30]) );
  NAND2X1 U1141 ( .A(n308), .B(n92), .Y(n54) );
  INVX2 U1142 ( .A(n91), .Y(n308) );
  OAI21X1 U1143 ( .A0(n101), .A1(n91), .B0(n92), .Y(n90) );
  INVX2 U1144 ( .A(n105), .Y(n103) );
  INVX2 U1145 ( .A(n116), .Y(n114) );
  NAND2X1 U1146 ( .A(n969), .B(n970), .Y(n100) );
  NOR2X1 U1147 ( .A(n100), .B(n91), .Y(n89) );
  ADDFX2 U1148 ( .A(n444), .B(n433), .CI(n431), .CO(n426), .S(n427) );
  ADDFHX1 U1149 ( .A(n485), .B(n483), .CI(n492), .CO(n478), .S(n479) );
  ADDFX2 U1150 ( .A(n529), .B(n532), .CI(n527), .CO(n524), .S(n525) );
  ADDFX2 U1151 ( .A(n535), .B(n538), .CI(n533), .CO(n530), .S(n531) );
  ADDFX2 U1152 ( .A(n513), .B(n518), .CI(n511), .CO(n508), .S(n509) );
  OR2X2 U1153 ( .A(n547), .B(n674), .Y(n965) );
  ADDFX2 U1154 ( .A(n514), .B(n512), .CI(n505), .CO(n500), .S(n501) );
  NAND2X1 U1155 ( .A(n691), .B(n563), .Y(n307) );
  NAND2X1 U1156 ( .A(n537), .B(n540), .Y(n288) );
  NOR2X1 U1157 ( .A(n690), .B(n675), .Y(n304) );
  OR2X1 U1158 ( .A(n541), .B(n544), .Y(n966) );
  OR2X1 U1159 ( .A(n537), .B(n540), .Y(n967) );
  AND2X1 U1160 ( .A(n944), .B(n307), .Y(product[1]) );
  NAND2X1 U1161 ( .A(n541), .B(n544), .Y(n294) );
  NAND2X1 U1162 ( .A(n545), .B(n546), .Y(n297) );
  NAND2XL U1163 ( .A(n690), .B(n675), .Y(n305) );
  NAND2X1 U1164 ( .A(n350), .B(n347), .Y(n140) );
  NAND2XL U1165 ( .A(n346), .B(n343), .Y(n129) );
  OR2X1 U1166 ( .A(n342), .B(n341), .Y(n969) );
  NAND2X1 U1167 ( .A(n342), .B(n341), .Y(n116) );
  INVX2 U1168 ( .A(n338), .Y(n339) );
  OR2X1 U1169 ( .A(n340), .B(n339), .Y(n970) );
  NAND2X1 U1170 ( .A(n340), .B(n339), .Y(n105) );
  NOR2X1 U1171 ( .A(n564), .B(n338), .Y(n91) );
  NAND2X1 U1172 ( .A(n564), .B(n338), .Y(n92) );
  OAI2BB1X1 U1173 ( .A0N(n867), .A1N(n6), .B0(n555), .Y(n676) );
  BUFX2 U1174 ( .A(n661), .Y(n971) );
  OAI22XL U1175 ( .A0(n30), .A1(n753), .B0(n752), .B1(n28), .Y(n618) );
  ADDFHX1 U1176 ( .A(n572), .B(n587), .CI(n602), .CO(n458), .S(n459) );
  OAI22XL U1177 ( .A0(n48), .A1(n707), .B0(n46), .B1(n706), .Y(n572) );
  ADDFHX1 U1178 ( .A(n646), .B(n586), .CI(n601), .CO(n444), .S(n445) );
  ADDFHX1 U1179 ( .A(n556), .B(n617), .CI(n632), .CO(n460), .S(n461) );
  OAI22XL U1180 ( .A0(n48), .A1(n868), .B0(n46), .B1(n708), .Y(n556) );
  OAI2BB1X1 U1181 ( .A0N(n9), .A1N(n12), .B0(n554), .Y(n659) );
  ADDFX2 U1182 ( .A(n613), .B(n643), .CI(n409), .CO(n406), .S(n407) );
  OAI2BB1X1 U1183 ( .A0N(n16), .A1N(n18), .B0(n553), .Y(n642) );
  INVX2 U1184 ( .A(n777), .Y(n553) );
  OAI2BB1X1 U1185 ( .A0N(n22), .A1N(n24), .B0(n552), .Y(n625) );
  INVX2 U1186 ( .A(n760), .Y(n552) );
  OAI22XL U1187 ( .A0(n42), .A1(n724), .B0(n723), .B1(n40), .Y(n589) );
  NOR2BXL U1188 ( .AN(b[0]), .B(n46), .Y(n573) );
  ADDFHX1 U1189 ( .A(n669), .B(n654), .CI(n534), .CO(n526), .S(n527) );
  ADDHXL U1190 ( .A(n685), .B(n655), .CO(n534), .S(n535) );
  ADDFHX1 U1191 ( .A(n560), .B(n640), .CI(n670), .CO(n532), .S(n533) );
  ADDFHX1 U1192 ( .A(n558), .B(n606), .CI(n666), .CO(n504), .S(n505) );
  ADDHXL U1193 ( .A(n683), .B(n653), .CO(n522), .S(n523) );
  ADDFHX1 U1194 ( .A(n668), .B(n523), .CI(n528), .CO(n518), .S(n519) );
  ADDFHX1 U1195 ( .A(n650), .B(n506), .CI(n497), .CO(n492), .S(n493) );
  ADDFHX1 U1196 ( .A(n583), .B(n598), .CI(n628), .CO(n404), .S(n405) );
  OAI22XL U1197 ( .A0(n30), .A1(n758), .B0(n757), .B1(n28), .Y(n623) );
  ADDFX2 U1198 ( .A(n658), .B(n688), .CI(n673), .CO(n544), .S(n545) );
  NOR2BXL U1199 ( .AN(b[0]), .B(n16), .Y(n658) );
  XNOR2X1 U1200 ( .A(b[0]), .B(n976), .Y(n775) );
  CLKINVXL U1201 ( .A(n972), .Y(n387) );
  INVX2 U1202 ( .A(n974), .Y(n874) );
  ADDFHX1 U1203 ( .A(n637), .B(n652), .CI(n667), .CO(n512), .S(n513) );
  NOR2BXL U1204 ( .AN(b[0]), .B(n40), .Y(n590) );
  ADDFX1 U1205 ( .A(n568), .B(n595), .CI(n610), .CO(n374), .S(n375) );
  OAI22XL U1206 ( .A0(n6), .A1(n875), .B0(n827), .B1(n867), .Y(n563) );
  INVX2 U1207 ( .A(n973), .Y(n875) );
  NAND2BX1 U1208 ( .AN(b[0]), .B(n973), .Y(n827) );
  XNOR2X1 U1209 ( .A(b[0]), .B(n979), .Y(n724) );
  ADDFHX1 U1210 ( .A(n570), .B(n584), .CI(n644), .CO(n418), .S(n419) );
  OAI2BB1X1 U1211 ( .A0N(n34), .A1N(n36), .B0(n550), .Y(n591) );
  NAND2BX1 U1212 ( .AN(b[0]), .B(n977), .Y(n759) );
  OAI22XL U1213 ( .A0(n826), .A1(n6), .B0(n825), .B1(n867), .Y(n691) );
  XNOR2X1 U1214 ( .A(b[0]), .B(n973), .Y(n826) );
  NOR2BXL U1215 ( .AN(b[0]), .B(n34), .Y(n607) );
  ADDFX2 U1216 ( .A(n368), .B(n578), .CI(n608), .CO(n360), .S(n361) );
  OAI2BB1X1 U1217 ( .A0N(n28), .A1N(n30), .B0(n551), .Y(n608) );
  INVX2 U1218 ( .A(n743), .Y(n551) );
  INVX1 U1219 ( .A(n368), .Y(n369) );
  NOR2BXL U1220 ( .AN(b[0]), .B(n28), .Y(n624) );
  ADDFHX1 U1221 ( .A(n641), .B(n686), .CI(n656), .CO(n538), .S(n539) );
  ADDHXL U1222 ( .A(n687), .B(n657), .CO(n542), .S(n543) );
  XNOR2X1 U1223 ( .A(b[0]), .B(n975), .Y(n792) );
  NAND2BX1 U1224 ( .AN(b[0]), .B(n980), .Y(n708) );
  NAND2BXL U1225 ( .AN(b[0]), .B(n979), .Y(n725) );
  XNOR2X1 U1226 ( .A(b[0]), .B(n974), .Y(n809) );
  ADDFX2 U1227 ( .A(n575), .B(n345), .CI(n348), .CO(n342), .S(n343) );
  INVX2 U1228 ( .A(n344), .Y(n345) );
  NAND2BX1 U1229 ( .AN(b[0]), .B(n974), .Y(n810) );
  XNOR2X1 U1230 ( .A(b[0]), .B(n977), .Y(n758) );
  NOR2BXL U1231 ( .AN(b[0]), .B(n9), .Y(n675) );
  NAND2BX1 U1232 ( .AN(b[0]), .B(n975), .Y(n793) );
  INVX2 U1233 ( .A(n979), .Y(n869) );
  INVX2 U1234 ( .A(n976), .Y(n872) );
  INVX2 U1235 ( .A(n980), .Y(n868) );
  INVX2 U1236 ( .A(n978), .Y(n870) );
  INVX2 U1237 ( .A(n977), .Y(n871) );
  NOR2BXL U1238 ( .AN(b[0]), .B(n867), .Y(product[0]) );
  ADDFX2 U1239 ( .A(n344), .B(n565), .CI(n574), .CO(n340), .S(n341) );
  OAI2BB1X1 U1240 ( .A0N(n40), .A1N(n42), .B0(n549), .Y(n574) );
  INVX2 U1241 ( .A(n709), .Y(n549) );
  OAI2BB1X1 U1242 ( .A0N(n46), .A1N(n48), .B0(n548), .Y(n564) );
  INVX2 U1243 ( .A(n692), .Y(n548) );
  XOR2X1 U1244 ( .A(n974), .B(a[2]), .Y(n850) );
  XOR2X1 U1245 ( .A(n979), .B(a[12]), .Y(n845) );
  XNOR2X1 U1246 ( .A(n973), .B(b[15]), .Y(n811) );
  XOR2X1 U1247 ( .A(n975), .B(a[4]), .Y(n849) );
  XNOR2X1 U1248 ( .A(n973), .B(b[11]), .Y(n815) );
  XOR2X1 U1249 ( .A(n976), .B(a[6]), .Y(n848) );
  XNOR2X1 U1250 ( .A(n973), .B(b[13]), .Y(n813) );
  XNOR2X1 U1251 ( .A(n973), .B(b[14]), .Y(n812) );
  XOR2X1 U1252 ( .A(n978), .B(a[10]), .Y(n846) );
  XNOR2X1 U1253 ( .A(n973), .B(b[10]), .Y(n816) );
  XNOR2X1 U1254 ( .A(n973), .B(b[12]), .Y(n814) );
  XNOR2X1 U1255 ( .A(n973), .B(b[7]), .Y(n819) );
  XNOR2X1 U1256 ( .A(n973), .B(b[9]), .Y(n817) );
  XNOR2X1 U1257 ( .A(n973), .B(b[6]), .Y(n820) );
  XNOR2X1 U1258 ( .A(n973), .B(b[4]), .Y(n822) );
  XNOR2X1 U1259 ( .A(n973), .B(b[8]), .Y(n818) );
  XNOR2X1 U1260 ( .A(n974), .B(b[15]), .Y(n794) );
  XNOR2X1 U1261 ( .A(n973), .B(b[3]), .Y(n823) );
  XNOR2X1 U1262 ( .A(n974), .B(b[12]), .Y(n797) );
  XNOR2X1 U1263 ( .A(n979), .B(b[3]), .Y(n721) );
  XNOR2X1 U1264 ( .A(n974), .B(b[11]), .Y(n798) );
  XNOR2X1 U1265 ( .A(n979), .B(b[4]), .Y(n720) );
  XNOR2X1 U1266 ( .A(n975), .B(b[11]), .Y(n781) );
  XNOR2X1 U1267 ( .A(n973), .B(b[2]), .Y(n824) );
  XNOR2X1 U1268 ( .A(n974), .B(b[14]), .Y(n795) );
  XNOR2X1 U1269 ( .A(n975), .B(b[7]), .Y(n785) );
  XNOR2X1 U1270 ( .A(n975), .B(b[12]), .Y(n780) );
  XNOR2X1 U1271 ( .A(n973), .B(b[5]), .Y(n821) );
  XNOR2X1 U1272 ( .A(n975), .B(b[9]), .Y(n783) );
  XNOR2X1 U1273 ( .A(n979), .B(b[2]), .Y(n722) );
  XNOR2X1 U1274 ( .A(n977), .B(b[8]), .Y(n750) );
  XNOR2X1 U1275 ( .A(n980), .B(b[1]), .Y(n706) );
  XNOR2X1 U1276 ( .A(n973), .B(b[1]), .Y(n825) );
  XNOR2X1 U1277 ( .A(n977), .B(b[6]), .Y(n752) );
  XNOR2X1 U1278 ( .A(n977), .B(b[9]), .Y(n749) );
  XNOR2X1 U1279 ( .A(n975), .B(b[10]), .Y(n782) );
  XNOR2X1 U1280 ( .A(n976), .B(b[10]), .Y(n765) );
  XNOR2X1 U1281 ( .A(n975), .B(b[6]), .Y(n786) );
  XNOR2X1 U1282 ( .A(n975), .B(b[3]), .Y(n789) );
  XNOR2X1 U1283 ( .A(n975), .B(b[8]), .Y(n784) );
  XNOR2X1 U1284 ( .A(n977), .B(b[7]), .Y(n751) );
  XNOR2X1 U1285 ( .A(n980), .B(b[5]), .Y(n702) );
  XNOR2X1 U1286 ( .A(n974), .B(b[10]), .Y(n799) );
  XNOR2X1 U1287 ( .A(n978), .B(b[8]), .Y(n733) );
  XNOR2X1 U1288 ( .A(n977), .B(b[5]), .Y(n753) );
  XNOR2X1 U1289 ( .A(n978), .B(b[4]), .Y(n737) );
  XNOR2X1 U1290 ( .A(n976), .B(b[9]), .Y(n766) );
  XNOR2X1 U1291 ( .A(n977), .B(b[11]), .Y(n747) );
  XNOR2X1 U1292 ( .A(n976), .B(b[8]), .Y(n767) );
  XNOR2X1 U1293 ( .A(n979), .B(b[5]), .Y(n719) );
  XNOR2X1 U1294 ( .A(n975), .B(b[2]), .Y(n790) );
  XNOR2X1 U1295 ( .A(n975), .B(b[5]), .Y(n787) );
  XNOR2X1 U1296 ( .A(n974), .B(b[13]), .Y(n796) );
  XNOR2X1 U1297 ( .A(n979), .B(b[1]), .Y(n723) );
  XNOR2X1 U1298 ( .A(n975), .B(b[14]), .Y(n778) );
  XNOR2X1 U1299 ( .A(n978), .B(b[7]), .Y(n734) );
  XNOR2X1 U1300 ( .A(n978), .B(b[3]), .Y(n738) );
  XNOR2X1 U1301 ( .A(n975), .B(b[4]), .Y(n788) );
  XNOR2X1 U1302 ( .A(n977), .B(b[10]), .Y(n748) );
  XNOR2X1 U1303 ( .A(n976), .B(b[6]), .Y(n769) );
  XNOR2X1 U1304 ( .A(n976), .B(b[7]), .Y(n768) );
  XNOR2X1 U1305 ( .A(n974), .B(b[9]), .Y(n800) );
  XNOR2X1 U1306 ( .A(n979), .B(b[8]), .Y(n716) );
  XNOR2X1 U1307 ( .A(n978), .B(b[9]), .Y(n732) );
  XNOR2X1 U1308 ( .A(n979), .B(b[10]), .Y(n714) );
  XNOR2X1 U1309 ( .A(n979), .B(b[7]), .Y(n717) );
  XNOR2X1 U1310 ( .A(n977), .B(b[4]), .Y(n754) );
  XNOR2X1 U1311 ( .A(n976), .B(b[15]), .Y(n760) );
  XNOR2X1 U1312 ( .A(n975), .B(b[13]), .Y(n779) );
  XNOR2X1 U1313 ( .A(n977), .B(b[3]), .Y(n755) );
  XNOR2X1 U1314 ( .A(n976), .B(b[1]), .Y(n774) );
  XNOR2X1 U1315 ( .A(n976), .B(b[5]), .Y(n770) );
  XNOR2X1 U1316 ( .A(n976), .B(b[4]), .Y(n771) );
  XNOR2X1 U1317 ( .A(n974), .B(b[2]), .Y(n807) );
  XNOR2X1 U1318 ( .A(n978), .B(b[12]), .Y(n729) );
  XNOR2X1 U1319 ( .A(n978), .B(b[2]), .Y(n739) );
  XNOR2X1 U1320 ( .A(n979), .B(b[9]), .Y(n715) );
  XNOR2X1 U1321 ( .A(n974), .B(b[6]), .Y(n803) );
  XNOR2X1 U1322 ( .A(n979), .B(b[6]), .Y(n718) );
  XNOR2X1 U1323 ( .A(n977), .B(b[2]), .Y(n756) );
  XNOR2X1 U1324 ( .A(n978), .B(b[11]), .Y(n730) );
  XNOR2X1 U1325 ( .A(n976), .B(b[3]), .Y(n772) );
  XNOR2X1 U1326 ( .A(n976), .B(b[2]), .Y(n773) );
  XNOR2X1 U1327 ( .A(n978), .B(b[1]), .Y(n740) );
  XNOR2X1 U1328 ( .A(n974), .B(b[1]), .Y(n808) );
  XNOR2X1 U1329 ( .A(n978), .B(b[10]), .Y(n731) );
  XNOR2X1 U1330 ( .A(n974), .B(b[5]), .Y(n804) );
  XNOR2X1 U1331 ( .A(n976), .B(b[14]), .Y(n761) );
  XNOR2X1 U1332 ( .A(n974), .B(b[3]), .Y(n806) );
  XNOR2X1 U1333 ( .A(n975), .B(b[1]), .Y(n791) );
  XNOR2X1 U1334 ( .A(n978), .B(b[5]), .Y(n736) );
  XNOR2X1 U1335 ( .A(n977), .B(b[1]), .Y(n757) );
  XNOR2X1 U1336 ( .A(n974), .B(b[4]), .Y(n805) );
  XNOR2X1 U1337 ( .A(n978), .B(b[6]), .Y(n735) );
  XNOR2X1 U1338 ( .A(n979), .B(b[11]), .Y(n713) );
  XNOR2X1 U1339 ( .A(n978), .B(b[13]), .Y(n728) );
  XNOR2X1 U1340 ( .A(n974), .B(b[7]), .Y(n802) );
  XNOR2X1 U1341 ( .A(n976), .B(b[11]), .Y(n764) );
  XNOR2X1 U1342 ( .A(n976), .B(b[12]), .Y(n763) );
  XNOR2X1 U1343 ( .A(n974), .B(b[8]), .Y(n801) );
  XNOR2X1 U1344 ( .A(n977), .B(b[12]), .Y(n746) );
  XNOR2X1 U1345 ( .A(n977), .B(b[14]), .Y(n744) );
  XNOR2X1 U1346 ( .A(n976), .B(b[13]), .Y(n762) );
  XNOR2X1 U1347 ( .A(n979), .B(b[13]), .Y(n711) );
  XNOR2X1 U1348 ( .A(n977), .B(b[13]), .Y(n745) );
  XNOR2X1 U1349 ( .A(n979), .B(b[14]), .Y(n710) );
  XNOR2X1 U1350 ( .A(n979), .B(b[12]), .Y(n712) );
  XNOR2X1 U1351 ( .A(n978), .B(b[15]), .Y(n726) );
  XNOR2X1 U1352 ( .A(n978), .B(b[14]), .Y(n727) );
  XNOR2X1 U1353 ( .A(n979), .B(b[15]), .Y(n709) );
  OAI22XL U1354 ( .A0(n12), .A1(n796), .B0(n795), .B1(n9), .Y(n661) );
  OAI22XL U1355 ( .A0(n30), .A1(n752), .B0(n751), .B1(n28), .Y(n617) );
  BUFX2 U1356 ( .A(n386), .Y(n972) );
  OAI22XL U1357 ( .A0(n48), .A1(n701), .B0(n46), .B1(n700), .Y(n386) );
  OAI22X1 U1358 ( .A0(n48), .A1(n706), .B0(n46), .B1(n705), .Y(n571) );
  ADDFHX1 U1359 ( .A(n408), .B(n597), .CI(n642), .CO(n396), .S(n397) );
  INVX1 U1360 ( .A(n408), .Y(n409) );
  OAI22XL U1361 ( .A0(n48), .A1(n703), .B0(n46), .B1(n702), .Y(n408) );
  OR2X1 U1362 ( .A(n631), .B(n571), .Y(n448) );
  AOI21XL U1363 ( .A0(n51), .A1(n118), .B0(n119), .Y(n117) );
  AOI21X4 U1364 ( .A0(n209), .A1(n222), .B0(n210), .Y(n208) );
  NOR2X4 U1365 ( .A(n389), .B(n398), .Y(n199) );
  OAI22X2 U1366 ( .A0(n48), .A1(n705), .B0(n46), .B1(n704), .Y(n434) );
  XOR2X2 U1367 ( .A(n229), .B(n68), .Y(product[16]) );
  NOR2XL U1368 ( .A(n53), .B(n109), .Y(n107) );
  NOR2X4 U1369 ( .A(n437), .B(n450), .Y(n227) );
  OAI22X1 U1370 ( .A0(n18), .A1(n792), .B0(n791), .B1(n16), .Y(n657) );
  OAI21XL U1371 ( .A0(n196), .A1(n188), .B0(n191), .Y(n187) );
  AOI21X4 U1372 ( .A0(n325), .A1(n251), .B0(n244), .Y(n242) );
  INVX4 U1373 ( .A(n245), .Y(n325) );
  XNOR2X1 U1374 ( .A(b[0]), .B(n978), .Y(n741) );
  AOI21X4 U1375 ( .A0(n255), .A1(n236), .B0(n237), .Y(n235) );
  ADDHX1 U1376 ( .A(n689), .B(n562), .CO(n546), .S(n547) );
  OAI21X1 U1377 ( .A0(n304), .A1(n307), .B0(n305), .Y(n303) );
endmodule


module PE_DW_mult_tc_31 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n6, n9, n12, n16, n18, n22, n24, n28, n30, n34, n36, n40, n42, n46,
         n48, n51, n52, n53, n54, n55, n56, n58, n59, n60, n61, n63, n64, n66,
         n67, n68, n69, n70, n71, n72, n74, n75, n76, n79, n80, n82, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n103, n105, n106, n107, n108, n109, n110, n114, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n140, n141,
         n142, n143, n144, n145, n148, n149, n151, n154, n155, n156, n157,
         n158, n159, n160, n164, n166, n167, n168, n169, n170, n171, n173,
         n176, n177, n181, n182, n183, n184, n185, n186, n187, n188, n191,
         n192, n193, n194, n196, n199, n200, n201, n203, n204, n205, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n219, n220,
         n221, n222, n224, n227, n228, n229, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n244, n246, n247, n248,
         n249, n251, n254, n255, n256, n257, n259, n261, n262, n264, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n281, n283, n284, n286, n288, n289, n290, n292, n294,
         n295, n296, n297, n298, n300, n302, n303, n304, n305, n307, n308,
         n311, n313, n315, n316, n319, n320, n322, n323, n324, n326, n329,
         n330, n334, n336, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n844, n845,
         n846, n847, n848, n849, n850, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997;

  AOI21X1 U60 ( .A0(n123), .A1(n89), .B0(n90), .Y(n88) );
  AOI21X1 U72 ( .A0(n123), .A1(n98), .B0(n99), .Y(n97) );
  AOI21X1 U76 ( .A0(n114), .A1(n987), .B0(n103), .Y(n101) );
  AOI21X1 U88 ( .A0(n123), .A1(n986), .B0(n114), .Y(n110) );
  AOI21X1 U106 ( .A0(n126), .A1(n151), .B0(n127), .Y(n125) );
  AOI21X1 U132 ( .A0(n160), .A1(n313), .B0(n151), .Y(n145) );
  NOR2X2 U169 ( .A(n370), .B(n363), .Y(n170) );
  NOR2X2 U203 ( .A(n389), .B(n398), .Y(n199) );
  NAND2X4 U212 ( .A(n399), .B(n410), .Y(n205) );
  OAI21X4 U214 ( .A0(n207), .A1(n235), .B0(n208), .Y(n51) );
  AOI21X1 U224 ( .A0(n214), .A1(n234), .B0(n215), .Y(n213) );
  ADDFHX4 U378 ( .A(n361), .B(n359), .CI(n364), .CO(n356), .S(n357) );
  ADDFHX4 U381 ( .A(n367), .B(n365), .CI(n372), .CO(n362), .S(n363) );
  ADDFHX4 U385 ( .A(n382), .B(n373), .CI(n380), .CO(n370), .S(n371) );
  ADDFHX4 U388 ( .A(n988), .B(n580), .CI(n625), .CO(n376), .S(n377) );
  ADDFHX4 U389 ( .A(n392), .B(n390), .CI(n381), .CO(n378), .S(n379) );
  ADDFHX4 U394 ( .A(n402), .B(n400), .CI(n391), .CO(n388), .S(n389) );
  ADDFHX4 U399 ( .A(n403), .B(n412), .CI(n401), .CO(n398), .S(n399) );
  ADDFHX4 U400 ( .A(n418), .B(n416), .CI(n414), .CO(n400), .S(n401) );
  ADDFHX4 U408 ( .A(n629), .B(n614), .CI(n432), .CO(n416), .S(n417) );
  ADDFHX4 U450 ( .A(n503), .B(n510), .CI(n501), .CO(n498), .S(n499) );
  OAI22X1 U555 ( .A0(n36), .A1(n732), .B0(n731), .B1(n34), .Y(n597) );
  OAI22X1 U557 ( .A0(n36), .A1(n734), .B0(n733), .B1(n34), .Y(n599) );
  OAI22X1 U560 ( .A0(n36), .A1(n737), .B0(n736), .B1(n34), .Y(n602) );
  OAI22X1 U561 ( .A0(n36), .A1(n738), .B0(n737), .B1(n34), .Y(n603) );
  OAI22X1 U562 ( .A0(n36), .A1(n739), .B0(n738), .B1(n34), .Y(n604) );
  OAI22X1 U563 ( .A0(n36), .A1(n740), .B0(n739), .B1(n34), .Y(n605) );
  OAI22X1 U586 ( .A0(n30), .A1(n744), .B0(n743), .B1(n28), .Y(n609) );
  OAI22X1 U587 ( .A0(n30), .A1(n745), .B0(n744), .B1(n28), .Y(n610) );
  OAI22X1 U588 ( .A0(n30), .A1(n746), .B0(n745), .B1(n28), .Y(n611) );
  OAI22X1 U589 ( .A0(n30), .A1(n747), .B0(n746), .B1(n28), .Y(n612) );
  OAI22X1 U591 ( .A0(n30), .A1(n749), .B0(n748), .B1(n28), .Y(n614) );
  OAI22X1 U592 ( .A0(n30), .A1(n750), .B0(n749), .B1(n28), .Y(n615) );
  OAI22X1 U593 ( .A0(n30), .A1(n751), .B0(n750), .B1(n28), .Y(n616) );
  OAI22X1 U594 ( .A0(n30), .A1(n752), .B0(n751), .B1(n28), .Y(n617) );
  OAI22X1 U597 ( .A0(n30), .A1(n755), .B0(n754), .B1(n28), .Y(n620) );
  OAI22X1 U598 ( .A0(n30), .A1(n756), .B0(n755), .B1(n28), .Y(n621) );
  OAI22X1 U599 ( .A0(n30), .A1(n757), .B0(n756), .B1(n28), .Y(n622) );
  OAI22X1 U622 ( .A0(n24), .A1(n761), .B0(n760), .B1(n968), .Y(n626) );
  OAI22X1 U623 ( .A0(n24), .A1(n762), .B0(n761), .B1(n968), .Y(n627) );
  OAI22X1 U624 ( .A0(n24), .A1(n763), .B0(n762), .B1(n968), .Y(n628) );
  OAI22X1 U625 ( .A0(n24), .A1(n764), .B0(n763), .B1(n968), .Y(n629) );
  OAI22X1 U626 ( .A0(n24), .A1(n765), .B0(n764), .B1(n968), .Y(n630) );
  OAI22X1 U627 ( .A0(n24), .A1(n766), .B0(n765), .B1(n968), .Y(n631) );
  OAI22X1 U628 ( .A0(n24), .A1(n767), .B0(n766), .B1(n968), .Y(n632) );
  OAI22X1 U629 ( .A0(n24), .A1(n768), .B0(n767), .B1(n968), .Y(n633) );
  OAI22X1 U630 ( .A0(n24), .A1(n769), .B0(n768), .B1(n968), .Y(n634) );
  OAI22X1 U631 ( .A0(n24), .A1(n770), .B0(n769), .B1(n968), .Y(n635) );
  OAI22X1 U632 ( .A0(n24), .A1(n771), .B0(n770), .B1(n968), .Y(n636) );
  OAI22X1 U633 ( .A0(n24), .A1(n772), .B0(n771), .B1(n22), .Y(n637) );
  OAI22X1 U634 ( .A0(n24), .A1(n773), .B0(n772), .B1(n968), .Y(n638) );
  OAI22X1 U635 ( .A0(n24), .A1(n774), .B0(n773), .B1(n968), .Y(n639) );
  OAI22X1 U655 ( .A0(n18), .A1(n873), .B0(n959), .B1(n793), .Y(n561) );
  OAI22X1 U658 ( .A0(n18), .A1(n778), .B0(n777), .B1(n959), .Y(n643) );
  OAI22X1 U659 ( .A0(n18), .A1(n779), .B0(n778), .B1(n959), .Y(n644) );
  OAI22X1 U660 ( .A0(n18), .A1(n780), .B0(n779), .B1(n959), .Y(n645) );
  OAI22X1 U661 ( .A0(n18), .A1(n781), .B0(n780), .B1(n959), .Y(n646) );
  OAI22X1 U663 ( .A0(n18), .A1(n783), .B0(n782), .B1(n959), .Y(n648) );
  OAI22X1 U665 ( .A0(n18), .A1(n785), .B0(n784), .B1(n959), .Y(n650) );
  OAI22X1 U667 ( .A0(n18), .A1(n787), .B0(n786), .B1(n959), .Y(n652) );
  OAI22X1 U669 ( .A0(n18), .A1(n789), .B0(n788), .B1(n959), .Y(n654) );
  OAI22X1 U671 ( .A0(n18), .A1(n791), .B0(n790), .B1(n959), .Y(n656) );
  OAI22X1 U698 ( .A0(n12), .A1(n799), .B0(n798), .B1(n9), .Y(n664) );
  OAI22X1 U730 ( .A0(n6), .A1(n812), .B0(n811), .B1(n867), .Y(n677) );
  OAI22X1 U732 ( .A0(n6), .A1(n814), .B0(n813), .B1(n867), .Y(n679) );
  OAI22X1 U733 ( .A0(n6), .A1(n815), .B0(n814), .B1(n867), .Y(n680) );
  OAI22X1 U734 ( .A0(n6), .A1(n816), .B0(n815), .B1(n867), .Y(n681) );
  OAI22X1 U735 ( .A0(n6), .A1(n817), .B0(n816), .B1(n867), .Y(n682) );
  OAI22X1 U736 ( .A0(n6), .A1(n818), .B0(n817), .B1(n867), .Y(n683) );
  OAI22X1 U737 ( .A0(n6), .A1(n819), .B0(n818), .B1(n867), .Y(n684) );
  OAI22X1 U738 ( .A0(n6), .A1(n820), .B0(n819), .B1(n867), .Y(n685) );
  OAI22X1 U739 ( .A0(n6), .A1(n821), .B0(n820), .B1(n867), .Y(n686) );
  OAI22X1 U740 ( .A0(n6), .A1(n822), .B0(n821), .B1(n867), .Y(n687) );
  OAI22X1 U741 ( .A0(n6), .A1(n823), .B0(n822), .B1(n867), .Y(n688) );
  OAI22X1 U742 ( .A0(n6), .A1(n824), .B0(n823), .B1(n867), .Y(n689) );
  OAI22X1 U743 ( .A0(n6), .A1(n825), .B0(n824), .B1(n867), .Y(n690) );
  NAND2X4 U786 ( .A(n46), .B(n844), .Y(n48) );
  NAND2X4 U789 ( .A(n40), .B(n845), .Y(n42) );
  NAND2X4 U792 ( .A(n34), .B(n846), .Y(n36) );
  XNOR2X4 U794 ( .A(n994), .B(a[10]), .Y(n34) );
  NAND2X4 U795 ( .A(n28), .B(n847), .Y(n30) );
  XNOR2X4 U797 ( .A(n993), .B(a[8]), .Y(n28) );
  NAND2X4 U798 ( .A(n22), .B(n848), .Y(n24) );
  NAND2X4 U801 ( .A(n958), .B(n849), .Y(n18) );
  XNOR2X4 U803 ( .A(n991), .B(a[4]), .Y(n16) );
  NAND2X4 U804 ( .A(n9), .B(n850), .Y(n12) );
  XNOR2X4 U806 ( .A(n990), .B(a[2]), .Y(n9) );
  ADDFHX4 U812 ( .A(n441), .B(n452), .CI(n439), .CO(n436), .S(n437) );
  OAI22XL U813 ( .A0(n36), .A1(n728), .B0(n727), .B1(n34), .Y(n593) );
  OAI22XL U814 ( .A0(n36), .A1(n727), .B0(n726), .B1(n34), .Y(n592) );
  OAI22XL U815 ( .A0(n36), .A1(n729), .B0(n728), .B1(n34), .Y(n594) );
  OAI22XL U816 ( .A0(n36), .A1(n735), .B0(n734), .B1(n34), .Y(n600) );
  OAI22XL U817 ( .A0(n36), .A1(n736), .B0(n735), .B1(n34), .Y(n601) );
  ADDFHX1 U818 ( .A(n633), .B(n603), .CI(n486), .CO(n470), .S(n471) );
  OAI21XL U819 ( .A0(n242), .A1(n238), .B0(n239), .Y(n237) );
  AOI21X2 U820 ( .A0(n960), .A1(n251), .B0(n244), .Y(n242) );
  OAI22X1 U821 ( .A0(n30), .A1(n754), .B0(n753), .B1(n28), .Y(n619) );
  NOR2X4 U822 ( .A(n411), .B(n422), .Y(n211) );
  OAI22X2 U823 ( .A0(n18), .A1(n782), .B0(n781), .B1(n959), .Y(n647) );
  XOR2X2 U824 ( .A(n677), .B(n647), .Y(n463) );
  XOR2X2 U825 ( .A(n201), .B(n64), .Y(product[20]) );
  XNOR2XL U826 ( .A(n997), .B(b[14]), .Y(n693) );
  XNOR2XL U827 ( .A(n996), .B(b[14]), .Y(n710) );
  OAI22XL U828 ( .A0(n12), .A1(n806), .B0(n805), .B1(n9), .Y(n671) );
  OAI22XL U829 ( .A0(n12), .A1(n808), .B0(n807), .B1(n9), .Y(n673) );
  OAI22XL U830 ( .A0(n12), .A1(n803), .B0(n802), .B1(n9), .Y(n668) );
  OAI22XL U831 ( .A0(n12), .A1(n805), .B0(n804), .B1(n9), .Y(n670) );
  OAI22XL U832 ( .A0(n12), .A1(n801), .B0(n800), .B1(n9), .Y(n666) );
  OAI22XL U833 ( .A0(n12), .A1(n802), .B0(n801), .B1(n9), .Y(n667) );
  OAI22XL U834 ( .A0(n12), .A1(n797), .B0(n796), .B1(n9), .Y(n662) );
  OAI22XL U835 ( .A0(n12), .A1(n804), .B0(n803), .B1(n9), .Y(n669) );
  OAI22XL U836 ( .A0(n12), .A1(n807), .B0(n806), .B1(n9), .Y(n672) );
  OAI22XL U837 ( .A0(n12), .A1(n795), .B0(n794), .B1(n9), .Y(n660) );
  OAI22XL U838 ( .A0(n12), .A1(n796), .B0(n795), .B1(n9), .Y(n661) );
  OAI22XL U839 ( .A0(n12), .A1(n798), .B0(n797), .B1(n9), .Y(n663) );
  INVX2 U840 ( .A(n943), .Y(n462) );
  NAND2XL U841 ( .A(n677), .B(n647), .Y(n943) );
  ADDFHX1 U842 ( .A(n662), .B(n463), .CI(n474), .CO(n456), .S(n457) );
  NAND2XL U843 ( .A(n996), .B(a[14]), .Y(n946) );
  NAND2X2 U844 ( .A(n944), .B(n945), .Y(n947) );
  NAND2X4 U845 ( .A(n946), .B(n947), .Y(n46) );
  INVXL U846 ( .A(n996), .Y(n944) );
  INVX2 U847 ( .A(a[14]), .Y(n945) );
  BUFX12 U848 ( .A(a[13]), .Y(n996) );
  OAI22XL U849 ( .A0(n48), .A1(n699), .B0(n46), .B1(n698), .Y(n368) );
  OAI22XL U850 ( .A0(n48), .A1(n700), .B0(n46), .B1(n699), .Y(n568) );
  OAI22XL U851 ( .A0(n48), .A1(n697), .B0(n46), .B1(n696), .Y(n354) );
  OAI22XL U852 ( .A0(n48), .A1(n698), .B0(n46), .B1(n697), .Y(n567) );
  OAI22XL U853 ( .A0(n48), .A1(n695), .B0(n46), .B1(n694), .Y(n344) );
  OAI22XL U854 ( .A0(n48), .A1(n696), .B0(n46), .B1(n695), .Y(n566) );
  OAI22XL U855 ( .A0(n48), .A1(n694), .B0(n46), .B1(n693), .Y(n565) );
  OAI22XL U856 ( .A0(n48), .A1(n693), .B0(n46), .B1(n692), .Y(n338) );
  NOR2BX1 U857 ( .AN(b[0]), .B(n46), .Y(n573) );
  NOR2X1 U858 ( .A(n46), .B(n705), .Y(n955) );
  OR2X2 U859 ( .A(n48), .B(n868), .Y(n948) );
  OR2X1 U860 ( .A(n46), .B(n708), .Y(n949) );
  NAND2X4 U861 ( .A(n948), .B(n949), .Y(n556) );
  CLKINVXL U862 ( .A(n997), .Y(n868) );
  NAND2BXL U863 ( .AN(b[0]), .B(n997), .Y(n708) );
  ADDFHX2 U864 ( .A(n556), .B(n617), .CI(n632), .CO(n460), .S(n461) );
  NAND2X1 U865 ( .A(n995), .B(a[12]), .Y(n952) );
  NAND2X2 U866 ( .A(n950), .B(n951), .Y(n953) );
  NAND2X4 U867 ( .A(n952), .B(n953), .Y(n40) );
  INVX1 U868 ( .A(n995), .Y(n950) );
  INVX4 U869 ( .A(a[12]), .Y(n951) );
  BUFX12 U870 ( .A(a[11]), .Y(n995) );
  OAI22XL U871 ( .A0(n42), .A1(n710), .B0(n709), .B1(n40), .Y(n575) );
  OAI22XL U872 ( .A0(n42), .A1(n711), .B0(n710), .B1(n40), .Y(n576) );
  OAI22XL U873 ( .A0(n42), .A1(n713), .B0(n712), .B1(n40), .Y(n578) );
  OAI22XL U874 ( .A0(n42), .A1(n714), .B0(n713), .B1(n40), .Y(n579) );
  OAI22XL U875 ( .A0(n42), .A1(n715), .B0(n714), .B1(n40), .Y(n580) );
  OAI22XL U876 ( .A0(n42), .A1(n723), .B0(n722), .B1(n40), .Y(n588) );
  OAI22XL U877 ( .A0(n42), .A1(n722), .B0(n721), .B1(n40), .Y(n587) );
  OAI22XL U878 ( .A0(n42), .A1(n719), .B0(n718), .B1(n40), .Y(n584) );
  OAI22XL U879 ( .A0(n42), .A1(n718), .B0(n717), .B1(n40), .Y(n583) );
  OAI22XL U880 ( .A0(n42), .A1(n717), .B0(n716), .B1(n40), .Y(n582) );
  OAI22X4 U881 ( .A0(n42), .A1(n869), .B0(n40), .B1(n725), .Y(n557) );
  NOR2XL U882 ( .A(n48), .B(n706), .Y(n954) );
  OR2X2 U883 ( .A(n954), .B(n955), .Y(n571) );
  OR2X2 U884 ( .A(n6), .B(n813), .Y(n956) );
  OR2X2 U885 ( .A(n812), .B(n867), .Y(n957) );
  NAND2X4 U886 ( .A(n956), .B(n957), .Y(n678) );
  INVX12 U887 ( .A(a[0]), .Y(n867) );
  ADDFHX2 U888 ( .A(n573), .B(n678), .CI(n588), .CO(n474), .S(n475) );
  ADDFHX1 U889 ( .A(n635), .B(n665), .CI(n620), .CO(n494), .S(n495) );
  XOR2X4 U890 ( .A(n997), .B(a[14]), .Y(n844) );
  ADDFHX1 U891 ( .A(n558), .B(n606), .CI(n666), .CO(n504), .S(n505) );
  BUFX8 U892 ( .A(n16), .Y(n958) );
  BUFX3 U893 ( .A(n16), .Y(n959) );
  INVX3 U894 ( .A(n235), .Y(n234) );
  ADDFHX1 U895 ( .A(n619), .B(n589), .CI(n604), .CO(n482), .S(n483) );
  OAI22X1 U896 ( .A0(n36), .A1(n741), .B0(n740), .B1(n34), .Y(n606) );
  XNOR2XL U897 ( .A(b[0]), .B(n995), .Y(n741) );
  OAI22X2 U898 ( .A0(n18), .A1(n786), .B0(n785), .B1(n959), .Y(n651) );
  XNOR2X2 U899 ( .A(n992), .B(b[11]), .Y(n781) );
  OAI22X1 U900 ( .A0(n42), .A1(n724), .B0(n723), .B1(n40), .Y(n589) );
  OAI21X2 U901 ( .A0(n211), .A1(n219), .B0(n212), .Y(n210) );
  XNOR2X2 U902 ( .A(n990), .B(b[12]), .Y(n814) );
  AOI21XL U903 ( .A0(n51), .A1(n85), .B0(n86), .Y(product[31]) );
  AOI21XL U904 ( .A0(n51), .A1(n94), .B0(n95), .Y(n93) );
  AOI21XL U905 ( .A0(n51), .A1(n118), .B0(n119), .Y(n117) );
  AOI21XL U906 ( .A0(n51), .A1(n131), .B0(n132), .Y(n130) );
  AOI21XL U907 ( .A0(n51), .A1(n168), .B0(n169), .Y(n167) );
  AOI21XL U908 ( .A0(n51), .A1(n155), .B0(n156), .Y(n154) );
  AOI21XL U909 ( .A0(n51), .A1(n177), .B0(n977), .Y(n176) );
  AOI21XL U910 ( .A0(n51), .A1(n186), .B0(n187), .Y(n185) );
  AOI21XL U911 ( .A0(n51), .A1(n193), .B0(n194), .Y(n192) );
  INVX4 U912 ( .A(n51), .Y(n963) );
  ADDFHX1 U913 ( .A(n557), .B(n664), .CI(n634), .CO(n484), .S(n485) );
  OAI21X2 U914 ( .A0(n227), .A1(n233), .B0(n228), .Y(n222) );
  NOR2X2 U915 ( .A(n437), .B(n450), .Y(n227) );
  NOR2X2 U916 ( .A(n423), .B(n436), .Y(n216) );
  ADDFHX2 U917 ( .A(n427), .B(n438), .CI(n425), .CO(n422), .S(n423) );
  BUFX12 U918 ( .A(a[9]), .Y(n994) );
  INVX2 U919 ( .A(n255), .Y(n254) );
  NAND2X1 U920 ( .A(n370), .B(n363), .Y(n171) );
  XNOR2X2 U921 ( .A(n992), .B(a[6]), .Y(n22) );
  NOR2X1 U922 ( .A(n690), .B(n675), .Y(n304) );
  NAND2X1 U923 ( .A(n691), .B(n563), .Y(n307) );
  ADDFX2 U924 ( .A(n568), .B(n595), .CI(n610), .CO(n374), .S(n375) );
  XNOR2X1 U925 ( .A(n273), .B(n75), .Y(product[9]) );
  ADDFX2 U926 ( .A(n594), .B(n579), .CI(n369), .CO(n366), .S(n367) );
  NAND2X1 U927 ( .A(n324), .B(n239), .Y(n70) );
  ADDFHX1 U928 ( .A(n493), .B(n500), .CI(n491), .CO(n488), .S(n489) );
  NOR2X1 U929 ( .A(n356), .B(n351), .Y(n148) );
  NAND2X1 U930 ( .A(n159), .B(n135), .Y(n133) );
  ADDFX2 U931 ( .A(n360), .B(n353), .CI(n358), .CO(n350), .S(n351) );
  ADDFX2 U932 ( .A(n566), .B(n352), .CI(n349), .CO(n346), .S(n347) );
  AOI21X1 U933 ( .A0(n269), .A1(n277), .B0(n270), .Y(n268) );
  NAND2X2 U934 ( .A(n989), .B(n498), .Y(n249) );
  NAND2XL U935 ( .A(n477), .B(n488), .Y(n246) );
  XOR2X1 U936 ( .A(n176), .B(n61), .Y(product[23]) );
  NAND2X1 U937 ( .A(n356), .B(n351), .Y(n149) );
  NOR2X1 U938 ( .A(n350), .B(n347), .Y(n137) );
  XOR2X1 U939 ( .A(n220), .B(n67), .Y(product[17]) );
  XOR2X1 U940 ( .A(n229), .B(n68), .Y(product[16]) );
  NAND2XL U941 ( .A(n322), .B(n228), .Y(n68) );
  NOR2X1 U942 ( .A(n346), .B(n343), .Y(n128) );
  ADDFHX1 U943 ( .A(n415), .B(n424), .CI(n413), .CO(n410), .S(n411) );
  ADDHXL U944 ( .A(n689), .B(n562), .CO(n546), .S(n547) );
  OAI22X1 U945 ( .A0(n826), .A1(n6), .B0(n825), .B1(n867), .Y(n691) );
  OAI22X1 U946 ( .A0(n6), .A1(n875), .B0(n827), .B1(n867), .Y(n563) );
  CMPR32X1 U947 ( .A(n560), .B(n640), .C(n670), .CO(n532), .S(n533) );
  CMPR32X1 U948 ( .A(n624), .B(n684), .C(n639), .CO(n528), .S(n529) );
  NAND2X2 U949 ( .A(n965), .B(n966), .Y(n653) );
  XOR2X1 U950 ( .A(n975), .B(n303), .Y(product[3]) );
  ADDFX2 U951 ( .A(n596), .B(n626), .CI(n387), .CO(n384), .S(n385) );
  ADDFX2 U952 ( .A(n637), .B(n652), .CI(n667), .CO(n512), .S(n513) );
  ADDFX2 U953 ( .A(n607), .B(n682), .CI(n622), .CO(n514), .S(n515) );
  ADDFX2 U954 ( .A(n636), .B(n621), .CI(n507), .CO(n502), .S(n503) );
  ADDFX2 U955 ( .A(n618), .B(n663), .CI(n648), .CO(n472), .S(n473) );
  XOR2X1 U956 ( .A(n284), .B(n974), .Y(product[7]) );
  AOI21X1 U957 ( .A0(n289), .A1(n985), .B0(n286), .Y(n284) );
  ADDFX2 U958 ( .A(n609), .B(n376), .CI(n374), .CO(n364), .S(n365) );
  XNOR2X1 U959 ( .A(n247), .B(n71), .Y(product[13]) );
  XOR2X1 U960 ( .A(n262), .B(n971), .Y(product[11]) );
  AOI21X1 U961 ( .A0(n267), .A1(n980), .B0(n264), .Y(n262) );
  ADDFX2 U962 ( .A(n567), .B(n593), .CI(n366), .CO(n358), .S(n359) );
  ADDFX2 U963 ( .A(n368), .B(n578), .CI(n608), .CO(n360), .S(n361) );
  ADDFX2 U964 ( .A(n592), .B(n577), .CI(n355), .CO(n352), .S(n353) );
  ADDFX2 U965 ( .A(n627), .B(n406), .CI(n404), .CO(n392), .S(n393) );
  ADDFX2 U966 ( .A(n611), .B(n581), .CI(n396), .CO(n382), .S(n383) );
  ADDFX2 U967 ( .A(n384), .B(n377), .CI(n375), .CO(n372), .S(n373) );
  ADDFX2 U968 ( .A(n394), .B(n385), .CI(n383), .CO(n380), .S(n381) );
  ADDFX2 U969 ( .A(n395), .B(n397), .CI(n393), .CO(n390), .S(n391) );
  NOR2X1 U970 ( .A(n489), .B(n498), .Y(n248) );
  ADDFX2 U971 ( .A(n650), .B(n506), .CI(n497), .CO(n492), .S(n493) );
  ADDFHX1 U972 ( .A(n514), .B(n512), .CI(n505), .CO(n500), .S(n501) );
  ADDFX2 U973 ( .A(n487), .B(n496), .CI(n494), .CO(n480), .S(n481) );
  ADDFHX1 U974 ( .A(n504), .B(n502), .CI(n495), .CO(n490), .S(n491) );
  ADDFX2 U975 ( .A(n572), .B(n587), .CI(n602), .CO(n458), .S(n459) );
  ADDFX2 U976 ( .A(n434), .B(n599), .CI(n659), .CO(n420), .S(n421) );
  ADDFX2 U977 ( .A(n646), .B(n586), .CI(n601), .CO(n444), .S(n445) );
  ADDFX2 U978 ( .A(n645), .B(n585), .CI(n630), .CO(n430), .S(n431) );
  ADDFX2 U979 ( .A(n615), .B(n660), .CI(n435), .CO(n432), .S(n433) );
  ADDFX2 U980 ( .A(n462), .B(n449), .CI(n460), .CO(n442), .S(n443) );
  XNOR2X1 U981 ( .A(n631), .B(n571), .Y(n449) );
  ADDFX2 U982 ( .A(n600), .B(n448), .CI(n446), .CO(n428), .S(n429) );
  OR2X1 U983 ( .A(n631), .B(n571), .Y(n448) );
  ADDFX2 U984 ( .A(n485), .B(n483), .CI(n492), .CO(n478), .S(n479) );
  ADDFX2 U985 ( .A(n475), .B(n484), .CI(n473), .CO(n468), .S(n469) );
  ADDFX2 U986 ( .A(n482), .B(n471), .CI(n480), .CO(n466), .S(n467) );
  ADDFX2 U987 ( .A(n472), .B(n470), .CI(n459), .CO(n454), .S(n455) );
  NOR2X1 U988 ( .A(n148), .B(n137), .Y(n135) );
  XNOR2X1 U989 ( .A(n234), .B(n69), .Y(product[15]) );
  BUFX8 U990 ( .A(a[15]), .Y(n997) );
  ADDFHX1 U991 ( .A(n481), .B(n490), .CI(n479), .CO(n476), .S(n477) );
  ADDFX2 U992 ( .A(n461), .B(n457), .CI(n468), .CO(n452), .S(n453) );
  ADDFX2 U993 ( .A(n458), .B(n447), .CI(n445), .CO(n440), .S(n441) );
  ADDFHX1 U994 ( .A(n428), .B(n417), .CI(n426), .CO(n412), .S(n413) );
  ADDFHX1 U995 ( .A(n444), .B(n433), .CI(n431), .CO(n426), .S(n427) );
  ADDFX2 U996 ( .A(n456), .B(n443), .CI(n454), .CO(n438), .S(n439) );
  ADDFHX1 U997 ( .A(n442), .B(n429), .CI(n440), .CO(n424), .S(n425) );
  ADDFX2 U998 ( .A(n469), .B(n478), .CI(n467), .CO(n464), .S(n465) );
  ADDFX2 U999 ( .A(n455), .B(n466), .CI(n453), .CO(n450), .S(n451) );
  NOR2X1 U1000 ( .A(n137), .B(n128), .Y(n126) );
  OAI21X1 U1001 ( .A0(n268), .A1(n256), .B0(n257), .Y(n255) );
  NAND2X1 U1002 ( .A(n979), .B(n980), .Y(n256) );
  NOR2X1 U1003 ( .A(n465), .B(n476), .Y(n238) );
  INVX2 U1004 ( .A(n249), .Y(n251) );
  NAND2X1 U1005 ( .A(n465), .B(n476), .Y(n239) );
  NAND2X1 U1006 ( .A(n451), .B(n464), .Y(n233) );
  NAND2X1 U1007 ( .A(n437), .B(n450), .Y(n228) );
  XOR2X1 U1008 ( .A(n117), .B(n56), .Y(product[28]) );
  NOR2X1 U1009 ( .A(n53), .B(n120), .Y(n118) );
  XOR2X1 U1010 ( .A(n106), .B(n55), .Y(product[29]) );
  NOR2X1 U1011 ( .A(n53), .B(n109), .Y(n107) );
  XOR2X1 U1012 ( .A(n167), .B(n60), .Y(product[24]) );
  NOR2X1 U1013 ( .A(n53), .B(n170), .Y(n168) );
  XOR2X1 U1014 ( .A(n154), .B(n59), .Y(product[25]) );
  NOR2X1 U1015 ( .A(n53), .B(n157), .Y(n155) );
  XOR2X1 U1016 ( .A(n141), .B(n58), .Y(product[26]) );
  XNOR2X1 U1017 ( .A(n130), .B(n972), .Y(product[27]) );
  NOR2X1 U1018 ( .A(n964), .B(n203), .Y(n201) );
  XOR2X1 U1019 ( .A(n192), .B(n63), .Y(product[21]) );
  INVX2 U1020 ( .A(n182), .Y(n978) );
  OAI21X1 U1021 ( .A0(n183), .A1(n191), .B0(n184), .Y(n182) );
  NOR2X1 U1022 ( .A(n204), .B(n199), .Y(n193) );
  AOI21X2 U1023 ( .A0(n255), .A1(n236), .B0(n237), .Y(n235) );
  NOR2X1 U1024 ( .A(n241), .B(n238), .Y(n236) );
  NAND2X1 U1025 ( .A(n423), .B(n436), .Y(n219) );
  NAND2X1 U1026 ( .A(n411), .B(n422), .Y(n212) );
  NOR2X2 U1027 ( .A(n211), .B(n216), .Y(n209) );
  NAND2X1 U1028 ( .A(n193), .B(n181), .Y(n53) );
  OR2X2 U1029 ( .A(n477), .B(n488), .Y(n960) );
  INVX2 U1030 ( .A(n977), .Y(n52) );
  OAI2BB1X1 U1031 ( .A0N(n194), .A1N(n181), .B0(n978), .Y(n977) );
  OR2X1 U1032 ( .A(n691), .B(n563), .Y(n961) );
  AND2X1 U1033 ( .A(n961), .B(n307), .Y(product[1]) );
  NOR2X1 U1034 ( .A(n399), .B(n410), .Y(n204) );
  AOI21X1 U1035 ( .A0(n979), .A1(n264), .B0(n259), .Y(n257) );
  OAI22X1 U1036 ( .A0(n18), .A1(n792), .B0(n791), .B1(n959), .Y(n657) );
  NOR2X1 U1037 ( .A(n963), .B(n204), .Y(n964) );
  OR2X2 U1038 ( .A(n18), .B(n788), .Y(n965) );
  OR2X1 U1039 ( .A(n787), .B(n959), .Y(n966) );
  ADDHX2 U1040 ( .A(n683), .B(n653), .CO(n522), .S(n523) );
  NAND2X2 U1041 ( .A(n315), .B(n981), .Y(n157) );
  CLKINVX3 U1042 ( .A(n22), .Y(n967) );
  AOI21XL U1043 ( .A0(n234), .A1(n323), .B0(n231), .Y(n229) );
  OAI21X1 U1044 ( .A0(n254), .A1(n248), .B0(n249), .Y(n247) );
  OAI21X1 U1045 ( .A0(n298), .A1(n296), .B0(n297), .Y(n295) );
  AND2X1 U1046 ( .A(n984), .B(n302), .Y(n975) );
  XOR2XL U1047 ( .A(n80), .B(n298), .Y(product[4]) );
  CLKINVXL U1048 ( .A(n296), .Y(n334) );
  AOI21XL U1049 ( .A0(n234), .A1(n221), .B0(n222), .Y(n220) );
  CLKINVXL U1050 ( .A(n290), .Y(n289) );
  NAND2XL U1051 ( .A(n509), .B(n516), .Y(n266) );
  INVX8 U1052 ( .A(n967), .Y(n968) );
  OAI21X4 U1053 ( .A0(n199), .A1(n205), .B0(n200), .Y(n194) );
  NAND2X1 U1054 ( .A(n389), .B(n398), .Y(n200) );
  INVX2 U1055 ( .A(n170), .Y(n315) );
  NAND2X2 U1056 ( .A(n388), .B(n379), .Y(n191) );
  XNOR2XL U1057 ( .A(n79), .B(n295), .Y(product[5]) );
  XOR2XL U1058 ( .A(n82), .B(n307), .Y(product[2]) );
  NAND2XL U1059 ( .A(n336), .B(n305), .Y(n82) );
  CLKINVXL U1060 ( .A(n304), .Y(n336) );
  NAND2BXL U1061 ( .AN(b[0]), .B(n991), .Y(n810) );
  XOR2X4 U1062 ( .A(n990), .B(a[0]), .Y(n976) );
  NAND2BX1 U1063 ( .AN(n216), .B(n219), .Y(n67) );
  XNOR2X1 U1064 ( .A(n185), .B(n970), .Y(product[22]) );
  CLKINVXL U1065 ( .A(n148), .Y(n313) );
  AND2X1 U1066 ( .A(n311), .B(n129), .Y(n972) );
  OAI21XL U1067 ( .A0(n149), .A1(n137), .B0(n140), .Y(n136) );
  NAND2XL U1068 ( .A(n982), .B(n283), .Y(n974) );
  OR2X4 U1069 ( .A(n531), .B(n536), .Y(n982) );
  OAI22XL U1070 ( .A0(n12), .A1(n874), .B0(n9), .B1(n810), .Y(n562) );
  ADDFX1 U1071 ( .A(n570), .B(n584), .CI(n644), .CO(n418), .S(n419) );
  CMPR32X1 U1072 ( .A(n569), .B(n582), .C(n612), .CO(n394), .S(n395) );
  ADDHXL U1073 ( .A(n679), .B(n649), .CO(n486), .S(n487) );
  XOR2X2 U1074 ( .A(n993), .B(a[6]), .Y(n848) );
  BUFX20 U1075 ( .A(a[5]), .Y(n992) );
  BUFX20 U1076 ( .A(a[3]), .Y(n991) );
  BUFX20 U1077 ( .A(a[1]), .Y(n990) );
  XOR2X1 U1078 ( .A(n994), .B(a[8]), .Y(n847) );
  XOR2X1 U1079 ( .A(n995), .B(a[10]), .Y(n846) );
  NOR2X1 U1080 ( .A(n53), .B(n133), .Y(n131) );
  XOR2X1 U1081 ( .A(n51), .B(n969), .Y(product[19]) );
  AND2X1 U1082 ( .A(n319), .B(n205), .Y(n969) );
  XOR2X1 U1083 ( .A(n213), .B(n66), .Y(product[18]) );
  NAND2XL U1084 ( .A(n320), .B(n212), .Y(n66) );
  NAND2BX1 U1085 ( .AN(n199), .B(n200), .Y(n64) );
  CLKINVXL U1086 ( .A(n232), .Y(n323) );
  NAND2XL U1087 ( .A(n159), .B(n313), .Y(n144) );
  AND2X1 U1088 ( .A(n316), .B(n184), .Y(n970) );
  NAND2XL U1089 ( .A(n315), .B(n171), .Y(n61) );
  AOI21X4 U1090 ( .A0(n981), .A1(n173), .B0(n164), .Y(n158) );
  INVX3 U1091 ( .A(n171), .Y(n173) );
  NAND2BX1 U1092 ( .AN(n188), .B(n191), .Y(n63) );
  NAND2XL U1093 ( .A(n313), .B(n149), .Y(n59) );
  NAND2XL U1094 ( .A(n979), .B(n261), .Y(n971) );
  NAND2XL U1095 ( .A(n330), .B(n275), .Y(n76) );
  CLKINVXL U1096 ( .A(n274), .Y(n330) );
  CLKINVXL U1097 ( .A(n277), .Y(n276) );
  NAND2XL U1098 ( .A(n329), .B(n272), .Y(n75) );
  OAI21XL U1099 ( .A0(n276), .A1(n274), .B0(n275), .Y(n273) );
  CLKINVXL U1100 ( .A(n271), .Y(n329) );
  NAND2X1 U1101 ( .A(n313), .B(n126), .Y(n124) );
  AOI21X1 U1102 ( .A0(n160), .A1(n135), .B0(n136), .Y(n134) );
  OR2X4 U1103 ( .A(n509), .B(n516), .Y(n980) );
  NAND2XL U1104 ( .A(n499), .B(n508), .Y(n261) );
  XOR2X1 U1105 ( .A(n254), .B(n72), .Y(product[12]) );
  NAND2BX1 U1106 ( .AN(n137), .B(n140), .Y(n58) );
  XOR2X1 U1107 ( .A(n973), .B(n289), .Y(product[6]) );
  AND2X1 U1108 ( .A(n985), .B(n288), .Y(n973) );
  NAND2XL U1109 ( .A(n362), .B(n357), .Y(n166) );
  NAND2XL U1110 ( .A(n983), .B(n294), .Y(n79) );
  OAI21XL U1111 ( .A0(n158), .A1(n124), .B0(n125), .Y(n123) );
  NAND2X1 U1112 ( .A(n122), .B(n986), .Y(n109) );
  ADDFHX1 U1113 ( .A(n522), .B(n515), .CI(n520), .CO(n510), .S(n511) );
  NAND2XL U1114 ( .A(n531), .B(n536), .Y(n283) );
  ADDFX1 U1115 ( .A(n521), .B(n526), .CI(n519), .CO(n516), .S(n517) );
  NAND2XL U1116 ( .A(n545), .B(n546), .Y(n297) );
  ADDFHX1 U1117 ( .A(n613), .B(n643), .CI(n409), .CO(n406), .S(n407) );
  OAI22XL U1118 ( .A0(n30), .A1(n748), .B0(n747), .B1(n28), .Y(n613) );
  OAI22XL U1119 ( .A0(n42), .A1(n716), .B0(n715), .B1(n40), .Y(n581) );
  ADDFHX1 U1120 ( .A(n590), .B(n680), .CI(n605), .CO(n496), .S(n497) );
  NOR2BXL U1121 ( .AN(b[0]), .B(n968), .Y(n641) );
  ADDFHX1 U1122 ( .A(n641), .B(n686), .CI(n656), .CO(n538), .S(n539) );
  CLKINVXL U1123 ( .A(n794), .Y(n554) );
  CMPR32X1 U1124 ( .A(n671), .B(n542), .C(n539), .CO(n536), .S(n537) );
  OAI22XL U1125 ( .A0(n30), .A1(n871), .B0(n28), .B1(n759), .Y(n559) );
  OAI22XL U1126 ( .A0(n36), .A1(n733), .B0(n732), .B1(n34), .Y(n598) );
  XNOR2XL U1127 ( .A(b[0]), .B(n994), .Y(n758) );
  OAI22XL U1128 ( .A0(n42), .A1(n720), .B0(n719), .B1(n40), .Y(n585) );
  ADDHXL U1129 ( .A(n685), .B(n655), .CO(n534), .S(n535) );
  OAI22XL U1130 ( .A0(n18), .A1(n790), .B0(n789), .B1(n959), .Y(n655) );
  OAI22XL U1131 ( .A0(n36), .A1(n870), .B0(n34), .B1(n742), .Y(n558) );
  XNOR2XL U1132 ( .A(b[0]), .B(n993), .Y(n775) );
  OAI22XL U1133 ( .A0(n30), .A1(n753), .B0(n752), .B1(n28), .Y(n618) );
  OAI22XL U1134 ( .A0(n48), .A1(n702), .B0(n46), .B1(n701), .Y(n569) );
  OAI22XL U1135 ( .A0(n42), .A1(n721), .B0(n720), .B1(n40), .Y(n586) );
  CMPR32X1 U1136 ( .A(n561), .B(n672), .C(n543), .CO(n540), .S(n541) );
  OAI22XL U1137 ( .A0(n48), .A1(n704), .B0(n46), .B1(n703), .Y(n570) );
  OAI22XL U1138 ( .A0(n12), .A1(n800), .B0(n799), .B1(n9), .Y(n665) );
  CLKINVXL U1139 ( .A(n760), .Y(n552) );
  XNOR2XL U1140 ( .A(b[0]), .B(n996), .Y(n724) );
  NAND2BXL U1141 ( .AN(b[0]), .B(n994), .Y(n759) );
  ADDHXL U1142 ( .A(n681), .B(n651), .CO(n506), .S(n507) );
  XNOR2X1 U1143 ( .A(b[0]), .B(n997), .Y(n707) );
  OAI22XL U1144 ( .A0(n18), .A1(n784), .B0(n783), .B1(n959), .Y(n649) );
  OAI22XL U1145 ( .A0(n36), .A1(n731), .B0(n730), .B1(n34), .Y(n596) );
  INVX1 U1146 ( .A(n368), .Y(n369) );
  OAI22XL U1147 ( .A0(n36), .A1(n730), .B0(n729), .B1(n34), .Y(n595) );
  OAI22XL U1148 ( .A0(n12), .A1(n809), .B0(n808), .B1(n9), .Y(n674) );
  NOR2BXL U1149 ( .AN(b[0]), .B(n9), .Y(n675) );
  CLKINVXL U1150 ( .A(n743), .Y(n551) );
  NAND2BXL U1151 ( .AN(b[0]), .B(n993), .Y(n776) );
  NAND2BXL U1152 ( .AN(b[0]), .B(n996), .Y(n725) );
  NAND2BXL U1153 ( .AN(b[0]), .B(n995), .Y(n742) );
  CLKINVXL U1154 ( .A(n994), .Y(n871) );
  CLKINVXL U1155 ( .A(n811), .Y(n555) );
  CLKINVXL U1156 ( .A(n993), .Y(n872) );
  CLKINVXL U1157 ( .A(n996), .Y(n869) );
  INVXL U1158 ( .A(n354), .Y(n355) );
  OAI22XL U1159 ( .A0(n42), .A1(n712), .B0(n711), .B1(n40), .Y(n577) );
  CLKINVXL U1160 ( .A(n995), .Y(n870) );
  NAND2X4 U1161 ( .A(n976), .B(n867), .Y(n6) );
  XOR2X1 U1162 ( .A(n991), .B(a[2]), .Y(n850) );
  XNOR2X1 U1163 ( .A(n997), .B(b[6]), .Y(n701) );
  XNOR2X1 U1164 ( .A(n997), .B(b[7]), .Y(n700) );
  XNOR2X1 U1165 ( .A(n997), .B(b[8]), .Y(n699) );
  XNOR2X1 U1166 ( .A(n997), .B(b[9]), .Y(n698) );
  XNOR2X1 U1167 ( .A(n997), .B(b[10]), .Y(n697) );
  XNOR2X1 U1168 ( .A(n997), .B(b[11]), .Y(n696) );
  XNOR2X1 U1169 ( .A(n997), .B(b[12]), .Y(n695) );
  XNOR2X1 U1170 ( .A(n997), .B(b[13]), .Y(n694) );
  XNOR2X1 U1171 ( .A(n997), .B(b[15]), .Y(n692) );
  NOR2X1 U1172 ( .A(n53), .B(n144), .Y(n142) );
  INVX2 U1173 ( .A(n122), .Y(n120) );
  NOR2X1 U1174 ( .A(n53), .B(n96), .Y(n94) );
  OAI21X1 U1175 ( .A0(n52), .A1(n157), .B0(n158), .Y(n156) );
  CLKINVXL U1176 ( .A(n211), .Y(n320) );
  NOR2X1 U1177 ( .A(n157), .B(n124), .Y(n122) );
  NOR2X1 U1178 ( .A(n227), .B(n232), .Y(n221) );
  CLKINVXL U1179 ( .A(n227), .Y(n322) );
  INVX2 U1180 ( .A(n268), .Y(n267) );
  OAI21XL U1181 ( .A0(n224), .A1(n216), .B0(n219), .Y(n215) );
  CLKINVXL U1182 ( .A(n222), .Y(n224) );
  NAND2XL U1183 ( .A(n323), .B(n233), .Y(n69) );
  INVX2 U1184 ( .A(n157), .Y(n159) );
  NOR2BXL U1185 ( .AN(n221), .B(n216), .Y(n214) );
  CLKINVXL U1186 ( .A(n204), .Y(n319) );
  CLKINVXL U1187 ( .A(n233), .Y(n231) );
  CLKINVXL U1188 ( .A(n205), .Y(n203) );
  NAND2XL U1189 ( .A(n122), .B(n98), .Y(n96) );
  NOR2X1 U1190 ( .A(n188), .B(n183), .Y(n181) );
  CLKINVXL U1191 ( .A(n53), .Y(n177) );
  INVX2 U1192 ( .A(n261), .Y(n259) );
  OAI21X1 U1193 ( .A0(n271), .A1(n275), .B0(n272), .Y(n270) );
  NOR2X1 U1194 ( .A(n271), .B(n274), .Y(n269) );
  OAI21XL U1195 ( .A0(n52), .A1(n170), .B0(n171), .Y(n169) );
  NAND2X1 U1196 ( .A(n981), .B(n166), .Y(n60) );
  NAND2X1 U1197 ( .A(n960), .B(n326), .Y(n241) );
  INVX2 U1198 ( .A(n248), .Y(n326) );
  NOR2X1 U1199 ( .A(n451), .B(n464), .Y(n232) );
  OAI21X1 U1200 ( .A0(n254), .A1(n241), .B0(n242), .Y(n240) );
  CLKINVXL U1201 ( .A(n238), .Y(n324) );
  INVX2 U1202 ( .A(n266), .Y(n264) );
  XNOR2X2 U1203 ( .A(n267), .B(n74), .Y(product[10]) );
  NAND2X1 U1204 ( .A(n980), .B(n266), .Y(n74) );
  OAI21XL U1205 ( .A0(n52), .A1(n120), .B0(n121), .Y(n119) );
  INVX2 U1206 ( .A(n123), .Y(n121) );
  CLKINVXL U1207 ( .A(n183), .Y(n316) );
  XOR2X1 U1208 ( .A(n276), .B(n76), .Y(product[8]) );
  NOR2BXL U1209 ( .AN(n193), .B(n188), .Y(n186) );
  INVX2 U1210 ( .A(n166), .Y(n164) );
  OAI21XL U1211 ( .A0(n196), .A1(n188), .B0(n191), .Y(n187) );
  CLKINVXL U1212 ( .A(n194), .Y(n196) );
  INVX2 U1213 ( .A(n149), .Y(n151) );
  OAI21XL U1214 ( .A0(n52), .A1(n96), .B0(n97), .Y(n95) );
  INVX2 U1215 ( .A(n101), .Y(n99) );
  NOR2X1 U1216 ( .A(n53), .B(n87), .Y(n85) );
  OAI21XL U1217 ( .A0(n52), .A1(n87), .B0(n88), .Y(n86) );
  NAND2XL U1218 ( .A(n122), .B(n89), .Y(n87) );
  INVX2 U1219 ( .A(n100), .Y(n98) );
  CLKINVXL U1220 ( .A(n128), .Y(n311) );
  NAND2X1 U1221 ( .A(n987), .B(n105), .Y(n55) );
  OAI21X1 U1222 ( .A0(n278), .A1(n290), .B0(n279), .Y(n277) );
  NAND2X1 U1223 ( .A(n982), .B(n985), .Y(n278) );
  AOI21X1 U1224 ( .A0(n982), .A1(n286), .B0(n281), .Y(n279) );
  INVX2 U1225 ( .A(n283), .Y(n281) );
  INVX2 U1226 ( .A(n246), .Y(n244) );
  OR2X4 U1227 ( .A(n499), .B(n508), .Y(n979) );
  NOR2X1 U1228 ( .A(n525), .B(n530), .Y(n274) );
  NAND2X1 U1229 ( .A(n986), .B(n116), .Y(n56) );
  AOI21X1 U1230 ( .A0(n295), .A1(n983), .B0(n292), .Y(n290) );
  INVX2 U1231 ( .A(n294), .Y(n292) );
  NOR2X1 U1232 ( .A(n517), .B(n524), .Y(n271) );
  AOI21X1 U1233 ( .A0(n984), .A1(n303), .B0(n300), .Y(n298) );
  INVX2 U1234 ( .A(n302), .Y(n300) );
  OAI21X1 U1235 ( .A0(n304), .A1(n307), .B0(n305), .Y(n303) );
  NAND2XL U1236 ( .A(n960), .B(n246), .Y(n71) );
  OAI21XL U1237 ( .A0(n140), .A1(n128), .B0(n129), .Y(n127) );
  NAND2X1 U1238 ( .A(n334), .B(n297), .Y(n80) );
  NAND2XL U1239 ( .A(n326), .B(n249), .Y(n72) );
  OR2X4 U1240 ( .A(n362), .B(n357), .Y(n981) );
  NAND2X1 U1241 ( .A(n517), .B(n524), .Y(n272) );
  INVX2 U1242 ( .A(n288), .Y(n286) );
  NAND2X1 U1243 ( .A(n525), .B(n530), .Y(n275) );
  NAND2X1 U1244 ( .A(n378), .B(n371), .Y(n184) );
  XOR2X1 U1245 ( .A(n93), .B(n54), .Y(product[30]) );
  NAND2X1 U1246 ( .A(n308), .B(n92), .Y(n54) );
  INVX2 U1247 ( .A(n91), .Y(n308) );
  OAI21X1 U1248 ( .A0(n101), .A1(n91), .B0(n92), .Y(n90) );
  INVX2 U1249 ( .A(n105), .Y(n103) );
  INVX2 U1250 ( .A(n116), .Y(n114) );
  NAND2X1 U1251 ( .A(n986), .B(n987), .Y(n100) );
  NOR2X1 U1252 ( .A(n100), .B(n91), .Y(n89) );
  ADDFHX1 U1253 ( .A(n430), .B(n421), .CI(n419), .CO(n414), .S(n415) );
  ADDFX2 U1254 ( .A(n535), .B(n538), .CI(n533), .CO(n530), .S(n531) );
  ADDFX2 U1255 ( .A(n529), .B(n532), .CI(n527), .CO(n524), .S(n525) );
  ADDFX2 U1256 ( .A(n513), .B(n518), .CI(n511), .CO(n508), .S(n509) );
  ADDFHX1 U1257 ( .A(n420), .B(n405), .CI(n407), .CO(n402), .S(n403) );
  OR2X1 U1258 ( .A(n541), .B(n544), .Y(n983) );
  OR2X1 U1259 ( .A(n547), .B(n674), .Y(n984) );
  NAND2X1 U1260 ( .A(n547), .B(n674), .Y(n302) );
  NOR2X1 U1261 ( .A(n545), .B(n546), .Y(n296) );
  NAND2X1 U1262 ( .A(n541), .B(n544), .Y(n294) );
  OR2X1 U1263 ( .A(n537), .B(n540), .Y(n985) );
  NAND2X1 U1264 ( .A(n537), .B(n540), .Y(n288) );
  NAND2X1 U1265 ( .A(n690), .B(n675), .Y(n305) );
  NAND2X1 U1266 ( .A(n350), .B(n347), .Y(n140) );
  NAND2XL U1267 ( .A(n346), .B(n343), .Y(n129) );
  OR2X1 U1268 ( .A(n342), .B(n341), .Y(n986) );
  NAND2X1 U1269 ( .A(n342), .B(n341), .Y(n116) );
  INVX2 U1270 ( .A(n338), .Y(n339) );
  OR2X1 U1271 ( .A(n340), .B(n339), .Y(n987) );
  NAND2X1 U1272 ( .A(n340), .B(n339), .Y(n105) );
  NOR2X1 U1273 ( .A(n564), .B(n338), .Y(n91) );
  NAND2X1 U1274 ( .A(n564), .B(n338), .Y(n92) );
  ADDFX2 U1275 ( .A(n408), .B(n597), .CI(n642), .CO(n396), .S(n397) );
  OAI2BB1X1 U1276 ( .A0N(n959), .A1N(n18), .B0(n553), .Y(n642) );
  INVX2 U1277 ( .A(n777), .Y(n553) );
  OAI2BB1X1 U1278 ( .A0N(n9), .A1N(n12), .B0(n554), .Y(n659) );
  OAI22XL U1279 ( .A0(n48), .A1(n705), .B0(n46), .B1(n704), .Y(n434) );
  OAI22XL U1280 ( .A0(n48), .A1(n707), .B0(n46), .B1(n706), .Y(n572) );
  OAI22XL U1281 ( .A0(n24), .A1(n872), .B0(n968), .B1(n776), .Y(n560) );
  OAI22XL U1282 ( .A0(n24), .A1(n775), .B0(n774), .B1(n968), .Y(n640) );
  OAI2BB1X1 U1283 ( .A0N(n968), .A1N(n24), .B0(n552), .Y(n625) );
  ADDFHX1 U1284 ( .A(n616), .B(n661), .CI(n676), .CO(n446), .S(n447) );
  OAI2BB1X1 U1285 ( .A0N(n867), .A1N(n6), .B0(n555), .Y(n676) );
  ADDFHX1 U1286 ( .A(n583), .B(n598), .CI(n628), .CO(n404), .S(n405) );
  ADDFHX1 U1287 ( .A(n559), .B(n623), .CI(n638), .CO(n520), .S(n521) );
  OAI22XL U1288 ( .A0(n30), .A1(n758), .B0(n757), .B1(n28), .Y(n623) );
  XNOR2X1 U1289 ( .A(b[0]), .B(n990), .Y(n826) );
  INVX2 U1290 ( .A(n990), .Y(n875) );
  NAND2BX1 U1291 ( .AN(b[0]), .B(n990), .Y(n827) );
  ADDHXL U1292 ( .A(n687), .B(n657), .CO(n542), .S(n543) );
  XNOR2X1 U1293 ( .A(b[0]), .B(n992), .Y(n792) );
  INVX2 U1294 ( .A(n992), .Y(n873) );
  ADDFHX1 U1295 ( .A(n668), .B(n523), .CI(n528), .CO(n518), .S(n519) );
  CMPR32X1 U1296 ( .A(n669), .B(n654), .C(n534), .CO(n526), .S(n527) );
  NOR2BXL U1297 ( .AN(b[0]), .B(n40), .Y(n590) );
  INVX2 U1298 ( .A(n991), .Y(n874) );
  ADDFX2 U1299 ( .A(n354), .B(n576), .CI(n591), .CO(n348), .S(n349) );
  OAI2BB1X1 U1300 ( .A0N(n34), .A1N(n36), .B0(n550), .Y(n591) );
  INVX2 U1301 ( .A(n726), .Y(n550) );
  NOR2BXL U1302 ( .AN(b[0]), .B(n28), .Y(n624) );
  NOR2BXL U1303 ( .AN(b[0]), .B(n34), .Y(n607) );
  NAND2BX1 U1304 ( .AN(b[0]), .B(n992), .Y(n793) );
  ADDFX2 U1305 ( .A(n658), .B(n688), .CI(n673), .CO(n544), .S(n545) );
  NOR2BX1 U1306 ( .AN(b[0]), .B(n959), .Y(n658) );
  CLKINVXL U1307 ( .A(n988), .Y(n387) );
  ADDFX2 U1308 ( .A(n575), .B(n345), .CI(n348), .CO(n342), .S(n343) );
  INVX2 U1309 ( .A(n344), .Y(n345) );
  OAI2BB1X1 U1310 ( .A0N(n28), .A1N(n30), .B0(n551), .Y(n608) );
  NOR2BXL U1311 ( .AN(b[0]), .B(n867), .Y(product[0]) );
  ADDFX2 U1312 ( .A(n344), .B(n565), .CI(n574), .CO(n340), .S(n341) );
  OAI2BB1X1 U1313 ( .A0N(n40), .A1N(n42), .B0(n549), .Y(n574) );
  INVX2 U1314 ( .A(n709), .Y(n549) );
  OAI2BB1X1 U1315 ( .A0N(n46), .A1N(n48), .B0(n548), .Y(n564) );
  INVX2 U1316 ( .A(n692), .Y(n548) );
  BUFX20 U1317 ( .A(a[7]), .Y(n993) );
  XOR2X1 U1318 ( .A(n992), .B(a[4]), .Y(n849) );
  XOR2X1 U1319 ( .A(n996), .B(a[12]), .Y(n845) );
  XNOR2X1 U1320 ( .A(n990), .B(b[15]), .Y(n811) );
  XNOR2X1 U1321 ( .A(n990), .B(b[11]), .Y(n815) );
  XNOR2X1 U1322 ( .A(n990), .B(b[13]), .Y(n813) );
  XNOR2X1 U1323 ( .A(n990), .B(b[10]), .Y(n816) );
  XNOR2X1 U1324 ( .A(n990), .B(b[9]), .Y(n817) );
  XNOR2X1 U1325 ( .A(n990), .B(b[7]), .Y(n819) );
  XNOR2X1 U1326 ( .A(n990), .B(b[14]), .Y(n812) );
  XNOR2X1 U1327 ( .A(n990), .B(b[8]), .Y(n818) );
  XNOR2X1 U1328 ( .A(n990), .B(b[6]), .Y(n820) );
  XNOR2X1 U1329 ( .A(n990), .B(b[4]), .Y(n822) );
  XNOR2X1 U1330 ( .A(n991), .B(b[15]), .Y(n794) );
  XNOR2X1 U1331 ( .A(n993), .B(b[10]), .Y(n765) );
  XNOR2X1 U1332 ( .A(n997), .B(b[5]), .Y(n702) );
  XNOR2X1 U1333 ( .A(n990), .B(b[3]), .Y(n823) );
  XNOR2X1 U1334 ( .A(n992), .B(b[15]), .Y(n777) );
  XNOR2X1 U1335 ( .A(n997), .B(b[3]), .Y(n704) );
  XNOR2X1 U1336 ( .A(n995), .B(b[8]), .Y(n733) );
  XNOR2X1 U1337 ( .A(n993), .B(b[9]), .Y(n766) );
  XNOR2X1 U1338 ( .A(n991), .B(b[12]), .Y(n797) );
  XNOR2X1 U1339 ( .A(n990), .B(b[1]), .Y(n825) );
  XNOR2X1 U1340 ( .A(n992), .B(b[7]), .Y(n785) );
  XNOR2X1 U1341 ( .A(n994), .B(b[6]), .Y(n752) );
  XNOR2X1 U1342 ( .A(n991), .B(b[14]), .Y(n795) );
  XNOR2X1 U1343 ( .A(n990), .B(b[2]), .Y(n824) );
  XNOR2X1 U1344 ( .A(n992), .B(b[9]), .Y(n783) );
  XNOR2X1 U1345 ( .A(n997), .B(b[4]), .Y(n703) );
  XNOR2X1 U1346 ( .A(n994), .B(b[9]), .Y(n749) );
  XNOR2X1 U1347 ( .A(n996), .B(b[4]), .Y(n720) );
  XNOR2X1 U1348 ( .A(n992), .B(b[10]), .Y(n782) );
  XNOR2X1 U1349 ( .A(n994), .B(b[11]), .Y(n747) );
  XNOR2X1 U1350 ( .A(n995), .B(b[7]), .Y(n734) );
  XNOR2X1 U1351 ( .A(n997), .B(b[2]), .Y(n705) );
  XNOR2X1 U1352 ( .A(n992), .B(b[12]), .Y(n780) );
  XNOR2X1 U1353 ( .A(n996), .B(b[5]), .Y(n719) );
  XNOR2X1 U1354 ( .A(n991), .B(b[11]), .Y(n798) );
  XNOR2X1 U1355 ( .A(n994), .B(b[8]), .Y(n750) );
  XNOR2X1 U1356 ( .A(n992), .B(b[6]), .Y(n786) );
  XNOR2X1 U1357 ( .A(n992), .B(b[13]), .Y(n779) );
  XNOR2X1 U1358 ( .A(n994), .B(b[5]), .Y(n753) );
  XNOR2X1 U1359 ( .A(n994), .B(b[7]), .Y(n751) );
  XNOR2X1 U1360 ( .A(n992), .B(b[14]), .Y(n778) );
  XNOR2X1 U1361 ( .A(n992), .B(b[8]), .Y(n784) );
  XNOR2X1 U1362 ( .A(n992), .B(b[3]), .Y(n789) );
  XNOR2X1 U1363 ( .A(n995), .B(b[9]), .Y(n732) );
  XNOR2X1 U1364 ( .A(n996), .B(b[3]), .Y(n721) );
  XNOR2X1 U1365 ( .A(n992), .B(b[5]), .Y(n787) );
  XNOR2X1 U1366 ( .A(n991), .B(b[13]), .Y(n796) );
  XNOR2X1 U1367 ( .A(n994), .B(b[10]), .Y(n748) );
  XNOR2X1 U1368 ( .A(n996), .B(b[7]), .Y(n717) );
  XNOR2X1 U1369 ( .A(n997), .B(b[1]), .Y(n706) );
  XNOR2X1 U1370 ( .A(n990), .B(b[5]), .Y(n821) );
  XNOR2X1 U1371 ( .A(n993), .B(b[4]), .Y(n771) );
  XNOR2X1 U1372 ( .A(n991), .B(b[10]), .Y(n799) );
  XNOR2X1 U1373 ( .A(n996), .B(b[6]), .Y(n718) );
  XNOR2X1 U1374 ( .A(n996), .B(b[2]), .Y(n722) );
  XNOR2X1 U1375 ( .A(n992), .B(b[2]), .Y(n790) );
  XNOR2X1 U1376 ( .A(n992), .B(b[4]), .Y(n788) );
  XNOR2X1 U1377 ( .A(n995), .B(b[4]), .Y(n737) );
  XNOR2X1 U1378 ( .A(n993), .B(b[6]), .Y(n769) );
  XNOR2X1 U1379 ( .A(n993), .B(b[3]), .Y(n772) );
  XNOR2X1 U1380 ( .A(n991), .B(b[9]), .Y(n800) );
  XNOR2X1 U1381 ( .A(n993), .B(b[8]), .Y(n767) );
  XNOR2X1 U1382 ( .A(n996), .B(b[1]), .Y(n723) );
  XNOR2X1 U1383 ( .A(n995), .B(b[2]), .Y(n739) );
  XNOR2X1 U1384 ( .A(n995), .B(b[1]), .Y(n740) );
  XNOR2X1 U1385 ( .A(n995), .B(b[3]), .Y(n738) );
  XNOR2X1 U1386 ( .A(n994), .B(b[4]), .Y(n754) );
  XNOR2X1 U1387 ( .A(n994), .B(b[3]), .Y(n755) );
  XNOR2X1 U1388 ( .A(n993), .B(b[5]), .Y(n770) );
  XNOR2X1 U1389 ( .A(n993), .B(b[7]), .Y(n768) );
  XNOR2X1 U1390 ( .A(n996), .B(b[10]), .Y(n714) );
  XNOR2X1 U1391 ( .A(n991), .B(b[3]), .Y(n806) );
  XNOR2X1 U1392 ( .A(n996), .B(b[8]), .Y(n716) );
  XNOR2X1 U1393 ( .A(n993), .B(b[1]), .Y(n774) );
  XNOR2X1 U1394 ( .A(n995), .B(b[10]), .Y(n731) );
  XNOR2X1 U1395 ( .A(n994), .B(b[2]), .Y(n756) );
  XNOR2X1 U1396 ( .A(n993), .B(b[15]), .Y(n760) );
  XNOR2X1 U1397 ( .A(n991), .B(b[6]), .Y(n803) );
  XNOR2X1 U1398 ( .A(n991), .B(b[2]), .Y(n807) );
  XNOR2X1 U1399 ( .A(n996), .B(b[9]), .Y(n715) );
  XNOR2X1 U1400 ( .A(n994), .B(b[1]), .Y(n757) );
  XNOR2X1 U1401 ( .A(n993), .B(b[2]), .Y(n773) );
  XNOR2X1 U1402 ( .A(n995), .B(b[11]), .Y(n730) );
  XNOR2X1 U1403 ( .A(n995), .B(b[12]), .Y(n729) );
  XNOR2X1 U1404 ( .A(n991), .B(b[1]), .Y(n808) );
  XNOR2X1 U1405 ( .A(n991), .B(b[5]), .Y(n804) );
  XNOR2X1 U1406 ( .A(n993), .B(b[14]), .Y(n761) );
  XNOR2X1 U1407 ( .A(n992), .B(b[1]), .Y(n791) );
  XNOR2X1 U1408 ( .A(n993), .B(b[12]), .Y(n763) );
  XNOR2X1 U1409 ( .A(n991), .B(b[8]), .Y(n801) );
  XNOR2X1 U1410 ( .A(n991), .B(b[4]), .Y(n805) );
  XNOR2X1 U1411 ( .A(n991), .B(b[7]), .Y(n802) );
  XNOR2X1 U1412 ( .A(n993), .B(b[11]), .Y(n764) );
  XNOR2X1 U1413 ( .A(n995), .B(b[6]), .Y(n735) );
  XNOR2X1 U1414 ( .A(n995), .B(b[5]), .Y(n736) );
  XNOR2X1 U1415 ( .A(n993), .B(b[13]), .Y(n762) );
  XNOR2X1 U1416 ( .A(n996), .B(b[11]), .Y(n713) );
  XNOR2X1 U1417 ( .A(n996), .B(b[13]), .Y(n711) );
  XNOR2X1 U1418 ( .A(n995), .B(b[13]), .Y(n728) );
  XNOR2X1 U1419 ( .A(n994), .B(b[12]), .Y(n746) );
  XNOR2X1 U1420 ( .A(n994), .B(b[13]), .Y(n745) );
  XNOR2X1 U1421 ( .A(n996), .B(b[12]), .Y(n712) );
  XNOR2X1 U1422 ( .A(n995), .B(b[15]), .Y(n726) );
  XNOR2X1 U1423 ( .A(n994), .B(b[14]), .Y(n744) );
  XNOR2X1 U1424 ( .A(n995), .B(b[14]), .Y(n727) );
  XNOR2X1 U1425 ( .A(n994), .B(b[15]), .Y(n743) );
  XNOR2X1 U1426 ( .A(n996), .B(b[15]), .Y(n709) );
  CLKINVXL U1427 ( .A(n434), .Y(n435) );
  XNOR2X1 U1428 ( .A(b[0]), .B(n991), .Y(n809) );
  BUFX2 U1429 ( .A(n386), .Y(n988) );
  OAI22XL U1430 ( .A0(n48), .A1(n701), .B0(n46), .B1(n700), .Y(n386) );
  INVX2 U1431 ( .A(n408), .Y(n409) );
  OAI22XL U1432 ( .A0(n48), .A1(n703), .B0(n46), .B1(n702), .Y(n408) );
  NAND2X2 U1433 ( .A(n209), .B(n221), .Y(n207) );
  XNOR2X2 U1434 ( .A(n240), .B(n70), .Y(product[14]) );
  AOI21X4 U1435 ( .A0(n209), .A1(n222), .B0(n210), .Y(n208) );
  XOR3X2 U1436 ( .A(n493), .B(n500), .C(n491), .Y(n989) );
  AOI21XL U1437 ( .A0(n51), .A1(n107), .B0(n108), .Y(n106) );
  OAI21X1 U1438 ( .A0(n52), .A1(n109), .B0(n110), .Y(n108) );
  OAI21XL U1439 ( .A0(n52), .A1(n144), .B0(n145), .Y(n143) );
  AOI21XL U1440 ( .A0(n51), .A1(n142), .B0(n143), .Y(n141) );
  NOR2X4 U1441 ( .A(n378), .B(n371), .Y(n183) );
  OAI21XL U1442 ( .A0(n52), .A1(n133), .B0(n134), .Y(n132) );
  INVX1 U1443 ( .A(n158), .Y(n160) );
  NOR2X4 U1444 ( .A(n388), .B(n379), .Y(n188) );
endmodule


module PE_DW_mult_tc_28 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n6, n9, n12, n16, n18, n22, n24, n28, n30, n34, n36, n40, n42, n46,
         n48, n51, n52, n53, n55, n56, n57, n58, n59, n61, n62, n63, n64, n66,
         n67, n68, n72, n73, n75, n76, n77, n80, n82, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n103,
         n105, n106, n107, n108, n109, n110, n114, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n140, n141, n142, n143,
         n144, n145, n148, n149, n151, n154, n155, n156, n157, n158, n159,
         n160, n164, n166, n167, n168, n169, n170, n171, n173, n176, n177,
         n181, n182, n183, n184, n185, n186, n187, n188, n191, n192, n193,
         n194, n196, n199, n200, n201, n203, n204, n205, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n219, n220, n221, n222,
         n224, n227, n228, n229, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n244, n246, n247, n248, n249, n251,
         n254, n255, n256, n257, n259, n261, n262, n264, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n281, n283, n284, n286, n288, n289, n290, n292, n294, n295, n296,
         n297, n298, n300, n302, n303, n304, n305, n307, n308, n313, n315,
         n316, n319, n320, n321, n323, n324, n326, n329, n330, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n844, n845, n846, n847, n848, n849, n850,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n943, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983;

  AOI21X1 U56 ( .A0(n972), .A1(n85), .B0(n86), .Y(product[31]) );
  AOI21X1 U60 ( .A0(n123), .A1(n89), .B0(n90), .Y(n88) );
  AOI21X1 U68 ( .A0(n972), .A1(n94), .B0(n95), .Y(n93) );
  AOI21X1 U72 ( .A0(n123), .A1(n98), .B0(n99), .Y(n97) );
  AOI21X1 U76 ( .A0(n114), .A1(n970), .B0(n103), .Y(n101) );
  AOI21X1 U84 ( .A0(n972), .A1(n107), .B0(n108), .Y(n106) );
  AOI21X1 U88 ( .A0(n123), .A1(n969), .B0(n114), .Y(n110) );
  AOI21X1 U106 ( .A0(n126), .A1(n151), .B0(n127), .Y(n125) );
  AOI21X1 U132 ( .A0(n160), .A1(n313), .B0(n151), .Y(n145) );
  AOI21X1 U144 ( .A0(n972), .A1(n155), .B0(n156), .Y(n154) );
  AOI21X1 U160 ( .A0(n972), .A1(n168), .B0(n169), .Y(n167) );
  AOI21X1 U172 ( .A0(n972), .A1(n177), .B0(n960), .Y(n176) );
  NOR2X2 U181 ( .A(n378), .B(n371), .Y(n183) );
  AOI21X1 U184 ( .A0(n972), .A1(n186), .B0(n187), .Y(n185) );
  NOR2X2 U191 ( .A(n388), .B(n379), .Y(n188) );
  NOR2X2 U203 ( .A(n389), .B(n398), .Y(n199) );
  NAND2X4 U212 ( .A(n399), .B(n410), .Y(n205) );
  NOR2X2 U239 ( .A(n227), .B(n232), .Y(n221) );
  NOR2X2 U251 ( .A(n451), .B(n464), .Y(n232) );
  NAND2X4 U252 ( .A(n451), .B(n464), .Y(n233) );
  AOI21X1 U255 ( .A0(n255), .A1(n236), .B0(n237), .Y(n235) );
  NAND2X4 U281 ( .A(n489), .B(n498), .Y(n249) );
  AOI21X1 U286 ( .A0(n946), .A1(n264), .B0(n259), .Y(n257) );
  ADDFHX4 U394 ( .A(n402), .B(n400), .CI(n391), .CO(n388), .S(n389) );
  ADDFHX4 U405 ( .A(n415), .B(n424), .CI(n413), .CO(n410), .S(n411) );
  ADDFHX4 U412 ( .A(n442), .B(n429), .CI(n440), .CO(n424), .S(n425) );
  ADDFHX4 U418 ( .A(n441), .B(n452), .CI(n439), .CO(n436), .S(n437) );
  ADDFHX4 U419 ( .A(n456), .B(n443), .CI(n454), .CO(n438), .S(n439) );
  ADDFHX4 U426 ( .A(n455), .B(n466), .CI(n453), .CO(n450), .S(n451) );
  ADDFHX4 U427 ( .A(n461), .B(n457), .CI(n468), .CO(n452), .S(n453) );
  ADDFHX4 U429 ( .A(n662), .B(n463), .CI(n474), .CO(n456), .S(n457) );
  ADDFHX4 U439 ( .A(n481), .B(n490), .CI(n479), .CO(n476), .S(n477) );
  ADDFHX4 U446 ( .A(n504), .B(n502), .CI(n495), .CO(n490), .S(n491) );
  ADDFHX4 U450 ( .A(n503), .B(n510), .CI(n501), .CO(n498), .S(n499) );
  OAI22X1 U475 ( .A0(n48), .A1(n868), .B0(n46), .B1(n708), .Y(n556) );
  OAI22X1 U478 ( .A0(n48), .A1(n693), .B0(n46), .B1(n692), .Y(n338) );
  OAI22X1 U479 ( .A0(n48), .A1(n694), .B0(n46), .B1(n693), .Y(n565) );
  OAI22X1 U480 ( .A0(n48), .A1(n695), .B0(n46), .B1(n694), .Y(n344) );
  OAI22X1 U481 ( .A0(n48), .A1(n696), .B0(n46), .B1(n695), .Y(n566) );
  OAI22X1 U482 ( .A0(n48), .A1(n697), .B0(n46), .B1(n696), .Y(n354) );
  OAI22X1 U483 ( .A0(n48), .A1(n698), .B0(n46), .B1(n697), .Y(n567) );
  OAI22X1 U484 ( .A0(n48), .A1(n699), .B0(n46), .B1(n698), .Y(n368) );
  OAI22X1 U485 ( .A0(n48), .A1(n700), .B0(n46), .B1(n699), .Y(n568) );
  OAI22X1 U486 ( .A0(n48), .A1(n701), .B0(n46), .B1(n700), .Y(n386) );
  OAI22X1 U487 ( .A0(n48), .A1(n702), .B0(n46), .B1(n701), .Y(n569) );
  OAI22X1 U488 ( .A0(n48), .A1(n703), .B0(n46), .B1(n702), .Y(n408) );
  OAI22X1 U489 ( .A0(n48), .A1(n704), .B0(n46), .B1(n703), .Y(n570) );
  OAI22X1 U491 ( .A0(n48), .A1(n706), .B0(n46), .B1(n705), .Y(n571) );
  OAI22X1 U511 ( .A0(n42), .A1(n869), .B0(n40), .B1(n725), .Y(n557) );
  OAI22X1 U514 ( .A0(n42), .A1(n710), .B0(n709), .B1(n40), .Y(n575) );
  OAI22X1 U515 ( .A0(n42), .A1(n711), .B0(n710), .B1(n40), .Y(n576) );
  OAI22X1 U517 ( .A0(n42), .A1(n713), .B0(n712), .B1(n40), .Y(n578) );
  OAI22X1 U519 ( .A0(n42), .A1(n715), .B0(n714), .B1(n40), .Y(n580) );
  OAI22X1 U522 ( .A0(n42), .A1(n718), .B0(n717), .B1(n40), .Y(n583) );
  OAI22X1 U527 ( .A0(n42), .A1(n723), .B0(n722), .B1(n40), .Y(n588) );
  OAI22X1 U528 ( .A0(n42), .A1(n724), .B0(n723), .B1(n40), .Y(n589) );
  OAI22X1 U547 ( .A0(n36), .A1(n870), .B0(n34), .B1(n742), .Y(n558) );
  OAI22X1 U550 ( .A0(n36), .A1(n727), .B0(n726), .B1(n34), .Y(n592) );
  OAI22X1 U551 ( .A0(n36), .A1(n728), .B0(n727), .B1(n34), .Y(n593) );
  OAI22X1 U552 ( .A0(n36), .A1(n729), .B0(n728), .B1(n34), .Y(n594) );
  OAI22X1 U554 ( .A0(n36), .A1(n731), .B0(n730), .B1(n34), .Y(n596) );
  OAI22X1 U555 ( .A0(n36), .A1(n732), .B0(n731), .B1(n34), .Y(n597) );
  OAI22X1 U557 ( .A0(n36), .A1(n734), .B0(n733), .B1(n34), .Y(n599) );
  OAI22X1 U559 ( .A0(n36), .A1(n736), .B0(n735), .B1(n34), .Y(n601) );
  OAI22X1 U560 ( .A0(n36), .A1(n737), .B0(n736), .B1(n34), .Y(n602) );
  OAI22X1 U561 ( .A0(n36), .A1(n738), .B0(n737), .B1(n34), .Y(n603) );
  OAI22X1 U562 ( .A0(n36), .A1(n739), .B0(n738), .B1(n34), .Y(n604) );
  OAI22X1 U563 ( .A0(n36), .A1(n740), .B0(n739), .B1(n34), .Y(n605) );
  OAI22X1 U564 ( .A0(n36), .A1(n741), .B0(n740), .B1(n34), .Y(n606) );
  OAI22X1 U583 ( .A0(n30), .A1(n871), .B0(n28), .B1(n759), .Y(n559) );
  OAI22X1 U586 ( .A0(n30), .A1(n744), .B0(n743), .B1(n28), .Y(n609) );
  OAI22X1 U587 ( .A0(n30), .A1(n745), .B0(n744), .B1(n28), .Y(n610) );
  OAI22X1 U588 ( .A0(n30), .A1(n746), .B0(n745), .B1(n28), .Y(n611) );
  OAI22X1 U589 ( .A0(n30), .A1(n747), .B0(n746), .B1(n28), .Y(n612) );
  OAI22X1 U590 ( .A0(n30), .A1(n748), .B0(n747), .B1(n28), .Y(n613) );
  OAI22X1 U591 ( .A0(n30), .A1(n749), .B0(n748), .B1(n28), .Y(n614) );
  OAI22X1 U592 ( .A0(n30), .A1(n750), .B0(n749), .B1(n28), .Y(n615) );
  OAI22X1 U596 ( .A0(n30), .A1(n754), .B0(n753), .B1(n28), .Y(n619) );
  OAI22X1 U597 ( .A0(n30), .A1(n755), .B0(n754), .B1(n28), .Y(n620) );
  OAI22X1 U598 ( .A0(n30), .A1(n756), .B0(n755), .B1(n28), .Y(n621) );
  OAI22X1 U599 ( .A0(n30), .A1(n757), .B0(n756), .B1(n28), .Y(n622) );
  OAI22X1 U619 ( .A0(n24), .A1(n872), .B0(n22), .B1(n776), .Y(n560) );
  OAI22X1 U623 ( .A0(n24), .A1(n762), .B0(n761), .B1(n22), .Y(n627) );
  OAI22X1 U624 ( .A0(n24), .A1(n763), .B0(n762), .B1(n22), .Y(n628) );
  OAI22X1 U625 ( .A0(n24), .A1(n764), .B0(n763), .B1(n22), .Y(n629) );
  OAI22X1 U626 ( .A0(n24), .A1(n765), .B0(n764), .B1(n22), .Y(n630) );
  OAI22X1 U627 ( .A0(n24), .A1(n766), .B0(n765), .B1(n22), .Y(n631) );
  OAI22X1 U628 ( .A0(n24), .A1(n767), .B0(n766), .B1(n22), .Y(n632) );
  OAI22X1 U629 ( .A0(n24), .A1(n768), .B0(n767), .B1(n22), .Y(n633) );
  OAI22X1 U630 ( .A0(n24), .A1(n769), .B0(n768), .B1(n22), .Y(n634) );
  OAI22X1 U632 ( .A0(n24), .A1(n771), .B0(n770), .B1(n22), .Y(n636) );
  OAI22X1 U633 ( .A0(n24), .A1(n772), .B0(n771), .B1(n22), .Y(n637) );
  OAI22X1 U634 ( .A0(n24), .A1(n773), .B0(n772), .B1(n22), .Y(n638) );
  OAI22X1 U635 ( .A0(n24), .A1(n774), .B0(n773), .B1(n22), .Y(n639) );
  OAI22X1 U655 ( .A0(n18), .A1(n873), .B0(n16), .B1(n793), .Y(n561) );
  OAI22X1 U659 ( .A0(n18), .A1(n779), .B0(n778), .B1(n16), .Y(n644) );
  OAI22X1 U660 ( .A0(n18), .A1(n780), .B0(n779), .B1(n16), .Y(n645) );
  OAI22X1 U661 ( .A0(n18), .A1(n781), .B0(n780), .B1(n16), .Y(n646) );
  OAI22X1 U662 ( .A0(n18), .A1(n782), .B0(n781), .B1(n16), .Y(n647) );
  OAI22X1 U663 ( .A0(n18), .A1(n783), .B0(n782), .B1(n16), .Y(n648) );
  OAI22X1 U665 ( .A0(n18), .A1(n785), .B0(n784), .B1(n16), .Y(n650) );
  OAI22X1 U667 ( .A0(n18), .A1(n787), .B0(n786), .B1(n16), .Y(n652) );
  OAI22X1 U671 ( .A0(n18), .A1(n791), .B0(n790), .B1(n16), .Y(n656) );
  OAI22X1 U672 ( .A0(n18), .A1(n792), .B0(n791), .B1(n16), .Y(n657) );
  OAI22X1 U694 ( .A0(n12), .A1(n795), .B0(n794), .B1(n9), .Y(n660) );
  OAI22X1 U696 ( .A0(n12), .A1(n797), .B0(n796), .B1(n9), .Y(n662) );
  OAI22X1 U697 ( .A0(n12), .A1(n798), .B0(n797), .B1(n9), .Y(n663) );
  OAI22X1 U699 ( .A0(n12), .A1(n800), .B0(n799), .B1(n9), .Y(n665) );
  OAI22X1 U700 ( .A0(n12), .A1(n801), .B0(n800), .B1(n9), .Y(n666) );
  OAI22X1 U701 ( .A0(n12), .A1(n802), .B0(n801), .B1(n9), .Y(n667) );
  OAI22X1 U702 ( .A0(n12), .A1(n803), .B0(n802), .B1(n9), .Y(n668) );
  OAI22X1 U703 ( .A0(n12), .A1(n804), .B0(n803), .B1(n9), .Y(n669) );
  OAI22X1 U704 ( .A0(n12), .A1(n805), .B0(n804), .B1(n9), .Y(n670) );
  OAI22X1 U705 ( .A0(n12), .A1(n806), .B0(n805), .B1(n9), .Y(n671) );
  OAI22X1 U706 ( .A0(n12), .A1(n807), .B0(n806), .B1(n9), .Y(n672) );
  OAI22X1 U707 ( .A0(n12), .A1(n808), .B0(n807), .B1(n9), .Y(n673) );
  OAI22X1 U708 ( .A0(n12), .A1(n809), .B0(n808), .B1(n9), .Y(n674) );
  OAI22X1 U727 ( .A0(n6), .A1(n875), .B0(n827), .B1(n867), .Y(n563) );
  OAI22X1 U730 ( .A0(n6), .A1(n812), .B0(n811), .B1(n867), .Y(n677) );
  OAI22X1 U731 ( .A0(n6), .A1(n813), .B0(n812), .B1(n867), .Y(n678) );
  OAI22X1 U732 ( .A0(n6), .A1(n814), .B0(n813), .B1(n867), .Y(n679) );
  OAI22X1 U733 ( .A0(n6), .A1(n815), .B0(n814), .B1(n867), .Y(n680) );
  OAI22X1 U734 ( .A0(n6), .A1(n816), .B0(n815), .B1(n867), .Y(n681) );
  OAI22X1 U735 ( .A0(n6), .A1(n817), .B0(n816), .B1(n867), .Y(n682) );
  OAI22X1 U736 ( .A0(n6), .A1(n818), .B0(n817), .B1(n867), .Y(n683) );
  OAI22X1 U737 ( .A0(n6), .A1(n819), .B0(n818), .B1(n867), .Y(n684) );
  OAI22X1 U738 ( .A0(n6), .A1(n820), .B0(n819), .B1(n867), .Y(n685) );
  OAI22X1 U739 ( .A0(n6), .A1(n821), .B0(n820), .B1(n867), .Y(n686) );
  OAI22X1 U740 ( .A0(n6), .A1(n822), .B0(n821), .B1(n867), .Y(n687) );
  OAI22X1 U741 ( .A0(n6), .A1(n823), .B0(n822), .B1(n867), .Y(n688) );
  OAI22X1 U742 ( .A0(n6), .A1(n824), .B0(n823), .B1(n867), .Y(n689) );
  OAI22X1 U743 ( .A0(n6), .A1(n825), .B0(n824), .B1(n867), .Y(n690) );
  OAI22X1 U744 ( .A0(n826), .A1(n6), .B0(n825), .B1(n867), .Y(n691) );
  NAND2X4 U786 ( .A(n46), .B(n844), .Y(n48) );
  XNOR2X4 U788 ( .A(n979), .B(a[14]), .Y(n46) );
  NAND2X4 U789 ( .A(n40), .B(n845), .Y(n42) );
  XNOR2X4 U791 ( .A(n978), .B(a[12]), .Y(n40) );
  NAND2X4 U792 ( .A(n34), .B(n846), .Y(n36) );
  XNOR2X4 U794 ( .A(n977), .B(a[10]), .Y(n34) );
  NAND2X4 U795 ( .A(n28), .B(n847), .Y(n30) );
  XNOR2X4 U797 ( .A(n976), .B(a[8]), .Y(n28) );
  NAND2X4 U798 ( .A(n22), .B(n848), .Y(n24) );
  XNOR2X4 U800 ( .A(n975), .B(a[6]), .Y(n22) );
  NAND2X4 U801 ( .A(n16), .B(n849), .Y(n18) );
  XNOR2X4 U803 ( .A(n974), .B(a[4]), .Y(n16) );
  NAND2X4 U804 ( .A(n9), .B(n850), .Y(n12) );
  XNOR2X4 U806 ( .A(n973), .B(a[2]), .Y(n9) );
  ADDHX1 U812 ( .A(n683), .B(n653), .CO(n522), .S(n523) );
  CLKINVX2 U813 ( .A(n277), .Y(n276) );
  OAI21X2 U814 ( .A0(n278), .A1(n290), .B0(n279), .Y(n277) );
  AOI21X4 U815 ( .A0(n965), .A1(n286), .B0(n281), .Y(n279) );
  AOI21X1 U816 ( .A0(n972), .A1(n193), .B0(n194), .Y(n192) );
  NOR2X2 U817 ( .A(n423), .B(n436), .Y(n216) );
  ADDFHX4 U818 ( .A(n427), .B(n438), .CI(n425), .CO(n422), .S(n423) );
  OAI21X2 U819 ( .A0(n207), .A1(n235), .B0(n208), .Y(n51) );
  AND2X4 U820 ( .A(n972), .B(n319), .Y(n943) );
  NOR2X4 U821 ( .A(n943), .B(n203), .Y(n201) );
  INVXL U822 ( .A(n204), .Y(n319) );
  CLKINVX12 U823 ( .A(n205), .Y(n203) );
  XOR2X4 U824 ( .A(n201), .B(n64), .Y(product[20]) );
  CMPR32X1 U825 ( .A(n434), .B(n599), .C(n659), .CO(n420), .S(n421) );
  OAI22X2 U826 ( .A0(n48), .A1(n705), .B0(n46), .B1(n704), .Y(n434) );
  ADDFHX1 U827 ( .A(n572), .B(n587), .CI(n602), .CO(n458), .S(n459) );
  OAI22XL U828 ( .A0(n48), .A1(n707), .B0(n46), .B1(n706), .Y(n572) );
  INVX1 U829 ( .A(n434), .Y(n435) );
  ADDFHX1 U830 ( .A(n556), .B(n617), .CI(n632), .CO(n460), .S(n461) );
  BUFX12 U831 ( .A(a[7]), .Y(n976) );
  BUFX12 U832 ( .A(a[9]), .Y(n977) );
  ADDFHX1 U833 ( .A(n616), .B(n661), .CI(n676), .CO(n446), .S(n447) );
  BUFX12 U834 ( .A(a[11]), .Y(n978) );
  ADDFHX1 U835 ( .A(n513), .B(n518), .CI(n511), .CO(n508), .S(n509) );
  NAND2X2 U836 ( .A(n509), .B(n516), .Y(n266) );
  ADDFHX1 U837 ( .A(n392), .B(n390), .CI(n381), .CO(n378), .S(n379) );
  ADDFX2 U838 ( .A(n566), .B(n352), .CI(n349), .CO(n346), .S(n347) );
  ADDFHX1 U839 ( .A(n382), .B(n373), .CI(n380), .CO(n370), .S(n371) );
  ADDFX2 U840 ( .A(n367), .B(n365), .CI(n372), .CO(n362), .S(n363) );
  NAND2X1 U841 ( .A(n370), .B(n363), .Y(n171) );
  NOR2X1 U842 ( .A(n399), .B(n410), .Y(n204) );
  NOR2X1 U843 ( .A(n346), .B(n343), .Y(n128) );
  NOR2X1 U844 ( .A(n370), .B(n363), .Y(n170) );
  ADDFHX1 U845 ( .A(n615), .B(n660), .CI(n435), .CO(n432), .S(n433) );
  ADDFHX1 U846 ( .A(n633), .B(n603), .CI(n486), .CO(n470), .S(n471) );
  ADDFX1 U847 ( .A(n613), .B(n643), .CI(n409), .CO(n406), .S(n407) );
  ADDFX2 U848 ( .A(n568), .B(n595), .CI(n610), .CO(n374), .S(n375) );
  XOR2X1 U849 ( .A(n973), .B(a[0]), .Y(n958) );
  ADDFHX1 U850 ( .A(n493), .B(n500), .CI(n491), .CO(n488), .S(n489) );
  ADDFX2 U851 ( .A(n594), .B(n579), .CI(n369), .CO(n366), .S(n367) );
  NOR2X1 U852 ( .A(n356), .B(n351), .Y(n148) );
  ADDFX2 U853 ( .A(n361), .B(n359), .CI(n364), .CO(n356), .S(n357) );
  ADDFX2 U854 ( .A(n360), .B(n353), .CI(n358), .CO(n350), .S(n351) );
  XOR2X1 U855 ( .A(n262), .B(n73), .Y(product[11]) );
  NOR2X1 U856 ( .A(n137), .B(n128), .Y(n126) );
  AOI21X1 U857 ( .A0(n963), .A1(n173), .B0(n164), .Y(n158) );
  INVX2 U858 ( .A(n171), .Y(n173) );
  NAND2X1 U859 ( .A(n313), .B(n126), .Y(n124) );
  NOR2X1 U860 ( .A(n350), .B(n347), .Y(n137) );
  OR2X2 U861 ( .A(n362), .B(n357), .Y(n963) );
  NAND2X1 U862 ( .A(n356), .B(n351), .Y(n149) );
  XOR2X1 U863 ( .A(n185), .B(n62), .Y(product[22]) );
  XOR2X1 U864 ( .A(n176), .B(n61), .Y(product[23]) );
  NAND2BXL U865 ( .AN(n199), .B(n200), .Y(n64) );
  XOR2X1 U866 ( .A(n130), .B(n57), .Y(product[27]) );
  NOR2X1 U867 ( .A(n53), .B(n133), .Y(n131) );
  NOR2X1 U868 ( .A(n53), .B(n120), .Y(n118) );
  NOR2X1 U869 ( .A(n53), .B(n109), .Y(n107) );
  NOR2X1 U870 ( .A(n53), .B(n96), .Y(n94) );
  NAND2X2 U871 ( .A(n193), .B(n181), .Y(n53) );
  NOR2X1 U872 ( .A(n12), .B(n799), .Y(n948) );
  NOR2X1 U873 ( .A(n798), .B(n9), .Y(n949) );
  ADDHXL U874 ( .A(n677), .B(n647), .CO(n462), .S(n463) );
  OAI22X1 U875 ( .A0(n18), .A1(n788), .B0(n787), .B1(n16), .Y(n653) );
  ADDFX2 U876 ( .A(n646), .B(n586), .CI(n601), .CO(n444), .S(n445) );
  ADDFX2 U877 ( .A(n637), .B(n652), .CI(n667), .CO(n512), .S(n513) );
  ADDFHX1 U878 ( .A(n514), .B(n512), .CI(n505), .CO(n500), .S(n501) );
  ADDFX2 U879 ( .A(n618), .B(n663), .CI(n648), .CO(n472), .S(n473) );
  ADDFX2 U880 ( .A(n573), .B(n678), .CI(n588), .CO(n474), .S(n475) );
  ADDHXL U881 ( .A(n679), .B(n649), .CO(n486), .S(n487) );
  ADDFX2 U882 ( .A(n635), .B(n665), .CI(n620), .CO(n494), .S(n495) );
  ADDFX2 U883 ( .A(n619), .B(n589), .CI(n604), .CO(n482), .S(n483) );
  ADDFHX1 U884 ( .A(n462), .B(n449), .CI(n460), .CO(n442), .S(n443) );
  XNOR2X1 U885 ( .A(n631), .B(n571), .Y(n449) );
  ADDFX2 U886 ( .A(n645), .B(n585), .CI(n630), .CO(n430), .S(n431) );
  ADDFX2 U887 ( .A(n600), .B(n448), .CI(n446), .CO(n428), .S(n429) );
  ADDFX2 U888 ( .A(n629), .B(n614), .CI(n432), .CO(n416), .S(n417) );
  ADDFX2 U889 ( .A(n570), .B(n584), .CI(n644), .CO(n418), .S(n419) );
  ADDFX2 U890 ( .A(n569), .B(n582), .CI(n612), .CO(n394), .S(n395) );
  ADDFX2 U891 ( .A(n596), .B(n626), .CI(n387), .CO(n384), .S(n385) );
  ADDHXL U892 ( .A(n689), .B(n562), .CO(n546), .S(n547) );
  ADDFX2 U893 ( .A(n658), .B(n688), .CI(n673), .CO(n544), .S(n545) );
  ADDFHX1 U894 ( .A(n472), .B(n470), .CI(n459), .CO(n454), .S(n455) );
  ADDFHX1 U895 ( .A(n458), .B(n447), .CI(n445), .CO(n440), .S(n441) );
  ADDFX2 U896 ( .A(n444), .B(n433), .CI(n431), .CO(n426), .S(n427) );
  ADDFX2 U897 ( .A(n482), .B(n471), .CI(n480), .CO(n466), .S(n467) );
  ADDFX2 U898 ( .A(n487), .B(n496), .CI(n494), .CO(n480), .S(n481) );
  ADDFX2 U899 ( .A(n430), .B(n421), .CI(n419), .CO(n414), .S(n415) );
  ADDFHX1 U900 ( .A(n428), .B(n417), .CI(n426), .CO(n412), .S(n413) );
  ADDFHX1 U901 ( .A(n418), .B(n416), .CI(n414), .CO(n400), .S(n401) );
  ADDFX2 U902 ( .A(n420), .B(n405), .CI(n407), .CO(n402), .S(n403) );
  ADDFX2 U903 ( .A(n627), .B(n406), .CI(n404), .CO(n392), .S(n393) );
  ADDFHX1 U904 ( .A(n395), .B(n397), .CI(n393), .CO(n390), .S(n391) );
  ADDFX2 U905 ( .A(n611), .B(n581), .CI(n396), .CO(n382), .S(n383) );
  ADDFX2 U906 ( .A(n394), .B(n385), .CI(n383), .CO(n380), .S(n381) );
  ADDFX2 U907 ( .A(n384), .B(n377), .CI(n375), .CO(n372), .S(n373) );
  ADDFX2 U908 ( .A(n609), .B(n376), .CI(n374), .CO(n364), .S(n365) );
  ADDFX2 U909 ( .A(n567), .B(n593), .CI(n366), .CO(n358), .S(n359) );
  ADDFX2 U910 ( .A(n368), .B(n578), .CI(n608), .CO(n360), .S(n361) );
  ADDFX2 U911 ( .A(n592), .B(n577), .CI(n355), .CO(n352), .S(n353) );
  NOR2X1 U912 ( .A(n545), .B(n546), .Y(n296) );
  NOR2X1 U913 ( .A(n489), .B(n498), .Y(n248) );
  BUFX8 U914 ( .A(a[13]), .Y(n979) );
  BUFX8 U915 ( .A(a[15]), .Y(n980) );
  ADDFHX1 U916 ( .A(n403), .B(n412), .CI(n401), .CO(n398), .S(n399) );
  NOR2X1 U917 ( .A(n148), .B(n137), .Y(n135) );
  NOR2X1 U918 ( .A(n690), .B(n675), .Y(n304) );
  NOR2X1 U919 ( .A(n411), .B(n422), .Y(n211) );
  OAI21X1 U920 ( .A0(n268), .A1(n256), .B0(n257), .Y(n255) );
  NOR2X1 U921 ( .A(n465), .B(n476), .Y(n238) );
  AOI21X2 U922 ( .A0(n947), .A1(n251), .B0(n244), .Y(n242) );
  INVX2 U923 ( .A(n249), .Y(n251) );
  AND2X1 U924 ( .A(n319), .B(n205), .Y(n959) );
  XOR2X1 U925 ( .A(n284), .B(n77), .Y(product[7]) );
  XOR2X1 U926 ( .A(n229), .B(n68), .Y(product[16]) );
  NAND2X1 U927 ( .A(n122), .B(n969), .Y(n109) );
  INVX2 U928 ( .A(n182), .Y(n961) );
  OAI21X1 U929 ( .A0(n183), .A1(n191), .B0(n184), .Y(n182) );
  OAI21X1 U930 ( .A0(n158), .A1(n124), .B0(n125), .Y(n123) );
  NOR2X1 U931 ( .A(n211), .B(n216), .Y(n209) );
  XOR2X1 U932 ( .A(n141), .B(n58), .Y(product[26]) );
  NOR2X1 U933 ( .A(n53), .B(n144), .Y(n142) );
  XNOR2X1 U934 ( .A(n167), .B(n953), .Y(product[24]) );
  NOR2X1 U935 ( .A(n53), .B(n170), .Y(n168) );
  XOR2X1 U936 ( .A(n154), .B(n59), .Y(product[25]) );
  NOR2X1 U937 ( .A(n53), .B(n157), .Y(n155) );
  INVX2 U938 ( .A(b[0]), .Y(n983) );
  INVX2 U939 ( .A(a[0]), .Y(n867) );
  XNOR2X1 U940 ( .A(n93), .B(n957), .Y(product[30]) );
  AND2X1 U941 ( .A(n966), .B(n307), .Y(product[1]) );
  INVX2 U942 ( .A(n960), .Y(n52) );
  OAI2BB1X1 U943 ( .A0N(n194), .A1N(n181), .B0(n961), .Y(n960) );
  OR2X2 U944 ( .A(n547), .B(n674), .Y(n945) );
  OR2X2 U945 ( .A(n499), .B(n508), .Y(n946) );
  OR2X2 U946 ( .A(n477), .B(n488), .Y(n947) );
  OAI22X1 U947 ( .A0(n12), .A1(n796), .B0(n795), .B1(n9), .Y(n661) );
  AOI21XL U948 ( .A0(n234), .A1(n221), .B0(n222), .Y(n220) );
  AOI21X1 U949 ( .A0(n209), .A1(n222), .B0(n210), .Y(n208) );
  XOR2X1 U950 ( .A(n192), .B(n63), .Y(product[21]) );
  OAI21X1 U951 ( .A0(n242), .A1(n238), .B0(n239), .Y(n237) );
  NAND2X1 U952 ( .A(n315), .B(n963), .Y(n157) );
  XOR2X1 U953 ( .A(n956), .B(n295), .Y(product[5]) );
  CLKINVXL U954 ( .A(n302), .Y(n300) );
  OR2X2 U955 ( .A(n948), .B(n949), .Y(n664) );
  NAND2BXL U956 ( .AN(n304), .B(n305), .Y(n82) );
  NOR2X1 U957 ( .A(n241), .B(n238), .Y(n236) );
  NOR2X1 U958 ( .A(n204), .B(n199), .Y(n193) );
  INVX1 U959 ( .A(n261), .Y(n259) );
  NAND2XL U960 ( .A(n946), .B(n964), .Y(n256) );
  NOR2BX1 U961 ( .AN(n193), .B(n188), .Y(n186) );
  INVX1 U962 ( .A(n288), .Y(n286) );
  CLKINVX2 U963 ( .A(n122), .Y(n120) );
  INVX2 U964 ( .A(n255), .Y(n254) );
  OAI21X1 U965 ( .A0(n199), .A1(n205), .B0(n200), .Y(n194) );
  NOR2X1 U966 ( .A(n525), .B(n530), .Y(n274) );
  INVX2 U967 ( .A(n148), .Y(n313) );
  NAND2X1 U968 ( .A(n477), .B(n488), .Y(n246) );
  INVX2 U969 ( .A(n235), .Y(n234) );
  AOI21XL U970 ( .A0(n234), .A1(n323), .B0(n231), .Y(n229) );
  NAND2XL U971 ( .A(n159), .B(n313), .Y(n144) );
  AOI21X1 U972 ( .A0(n269), .A1(n277), .B0(n270), .Y(n268) );
  XOR2X1 U973 ( .A(n972), .B(n959), .Y(product[19]) );
  NAND2BX1 U974 ( .AN(n188), .B(n191), .Y(n63) );
  OAI21X2 U975 ( .A0(n227), .A1(n233), .B0(n228), .Y(n222) );
  OAI21XL U976 ( .A0(n211), .A1(n219), .B0(n212), .Y(n210) );
  NAND2BXL U977 ( .AN(n227), .B(n228), .Y(n68) );
  AND2X1 U978 ( .A(n963), .B(n166), .Y(n953) );
  NOR2X2 U979 ( .A(n188), .B(n183), .Y(n181) );
  NAND2X1 U980 ( .A(n159), .B(n135), .Y(n133) );
  AOI21XL U981 ( .A0(n972), .A1(n131), .B0(n132), .Y(n130) );
  AOI21XL U982 ( .A0(n972), .A1(n142), .B0(n143), .Y(n141) );
  NAND2XL U983 ( .A(n965), .B(n283), .Y(n77) );
  NAND2XL U984 ( .A(n378), .B(n371), .Y(n184) );
  ADDFHX2 U985 ( .A(n521), .B(n526), .CI(n519), .CO(n516), .S(n517) );
  ADDFHX1 U986 ( .A(n485), .B(n483), .CI(n492), .CO(n478), .S(n479) );
  ADDFHX1 U987 ( .A(n522), .B(n515), .CI(n520), .CO(n510), .S(n511) );
  OR2X4 U988 ( .A(n531), .B(n536), .Y(n965) );
  INVX1 U989 ( .A(n408), .Y(n409) );
  ADDFX1 U990 ( .A(n669), .B(n654), .CI(n534), .CO(n526), .S(n527) );
  CMPR32X1 U991 ( .A(n671), .B(n542), .C(n539), .CO(n536), .S(n537) );
  OR2X1 U992 ( .A(n631), .B(n571), .Y(n448) );
  BUFX20 U993 ( .A(a[3]), .Y(n974) );
  XNOR2X1 U994 ( .A(n980), .B(b[5]), .Y(n702) );
  XNOR2X1 U995 ( .A(n980), .B(b[6]), .Y(n701) );
  XNOR2X1 U996 ( .A(n980), .B(b[10]), .Y(n697) );
  XNOR2X1 U997 ( .A(n980), .B(b[11]), .Y(n696) );
  XOR2X1 U998 ( .A(n240), .B(n950), .Y(product[14]) );
  AND2X1 U999 ( .A(n324), .B(n239), .Y(n950) );
  XOR2X1 U1000 ( .A(n234), .B(n951), .Y(product[15]) );
  AND2X1 U1001 ( .A(n323), .B(n233), .Y(n951) );
  XOR2X1 U1002 ( .A(n213), .B(n66), .Y(product[18]) );
  NAND2XL U1003 ( .A(n320), .B(n212), .Y(n66) );
  XOR2X1 U1004 ( .A(n220), .B(n67), .Y(product[17]) );
  NAND2XL U1005 ( .A(n321), .B(n219), .Y(n67) );
  OAI21XL U1006 ( .A0(n52), .A1(n144), .B0(n145), .Y(n143) );
  NAND2X1 U1007 ( .A(n437), .B(n450), .Y(n228) );
  XOR2X1 U1008 ( .A(n267), .B(n952), .Y(product[10]) );
  AND2X1 U1009 ( .A(n964), .B(n266), .Y(n952) );
  NAND2X1 U1010 ( .A(n947), .B(n326), .Y(n241) );
  AOI21XL U1011 ( .A0(n267), .A1(n964), .B0(n264), .Y(n262) );
  XOR2X1 U1012 ( .A(n247), .B(n954), .Y(product[13]) );
  AND2X1 U1013 ( .A(n947), .B(n246), .Y(n954) );
  NAND2XL U1014 ( .A(n313), .B(n149), .Y(n59) );
  XNOR2X1 U1015 ( .A(n273), .B(n75), .Y(product[9]) );
  OAI21X1 U1016 ( .A0(n276), .A1(n274), .B0(n275), .Y(n273) );
  CLKINVXL U1017 ( .A(n271), .Y(n329) );
  INVX2 U1018 ( .A(n170), .Y(n315) );
  NAND2XL U1019 ( .A(n499), .B(n508), .Y(n261) );
  NAND2BX1 U1020 ( .AN(n137), .B(n140), .Y(n58) );
  NAND2XL U1021 ( .A(n517), .B(n524), .Y(n272) );
  NAND2BX1 U1022 ( .AN(n128), .B(n129), .Y(n57) );
  NAND2XL U1023 ( .A(n525), .B(n530), .Y(n275) );
  XOR2X1 U1024 ( .A(n955), .B(n289), .Y(product[6]) );
  AND2X1 U1025 ( .A(n968), .B(n288), .Y(n955) );
  AOI21XL U1026 ( .A0(n289), .A1(n968), .B0(n286), .Y(n284) );
  AND2X1 U1027 ( .A(n967), .B(n294), .Y(n956) );
  XOR2XL U1028 ( .A(n962), .B(n303), .Y(product[3]) );
  OAI21XL U1029 ( .A0(n52), .A1(n133), .B0(n134), .Y(n132) );
  NAND2BX1 U1030 ( .AN(n296), .B(n297), .Y(n80) );
  NAND2XL U1031 ( .A(n362), .B(n357), .Y(n166) );
  AND2X1 U1032 ( .A(n308), .B(n92), .Y(n957) );
  NAND2XL U1033 ( .A(n531), .B(n536), .Y(n283) );
  NAND2XL U1034 ( .A(n545), .B(n546), .Y(n297) );
  ADDFHX1 U1035 ( .A(n557), .B(n664), .CI(n634), .CO(n484), .S(n485) );
  ADDFHX1 U1036 ( .A(n590), .B(n680), .CI(n605), .CO(n496), .S(n497) );
  ADDFHX1 U1037 ( .A(n641), .B(n686), .CI(n656), .CO(n538), .S(n539) );
  ADDFHX1 U1038 ( .A(n607), .B(n682), .CI(n622), .CO(n514), .S(n515) );
  CMPR32X1 U1039 ( .A(n668), .B(n523), .C(n528), .CO(n518), .S(n519) );
  ADDHXL U1040 ( .A(n681), .B(n651), .CO(n506), .S(n507) );
  OAI22XL U1041 ( .A0(n18), .A1(n786), .B0(n785), .B1(n16), .Y(n651) );
  OAI22XL U1042 ( .A0(n30), .A1(n753), .B0(n752), .B1(n28), .Y(n618) );
  OAI22XL U1043 ( .A0(n36), .A1(n735), .B0(n734), .B1(n34), .Y(n600) );
  OAI22XL U1044 ( .A0(n24), .A1(n770), .B0(n769), .B1(n22), .Y(n635) );
  OAI22XL U1045 ( .A0(n18), .A1(n789), .B0(n788), .B1(n16), .Y(n654) );
  OAI22XL U1046 ( .A0(n30), .A1(n752), .B0(n751), .B1(n28), .Y(n617) );
  OAI22XL U1047 ( .A0(n42), .A1(n721), .B0(n720), .B1(n40), .Y(n586) );
  OAI22XL U1048 ( .A0(n18), .A1(n790), .B0(n789), .B1(n16), .Y(n655) );
  OAI22XL U1049 ( .A0(n30), .A1(n758), .B0(n757), .B1(n28), .Y(n623) );
  OAI22XL U1050 ( .A0(n18), .A1(n784), .B0(n783), .B1(n16), .Y(n649) );
  OAI22XL U1051 ( .A0(n42), .A1(n720), .B0(n719), .B1(n40), .Y(n585) );
  OAI22XL U1052 ( .A0(n30), .A1(n751), .B0(n750), .B1(n28), .Y(n616) );
  OAI22XL U1053 ( .A0(n42), .A1(n716), .B0(n715), .B1(n40), .Y(n581) );
  CLKINVXL U1054 ( .A(n975), .Y(n873) );
  ADDFX1 U1055 ( .A(n561), .B(n672), .CI(n543), .CO(n540), .S(n541) );
  OAI22XL U1056 ( .A0(n18), .A1(n778), .B0(n777), .B1(n16), .Y(n643) );
  XNOR2XL U1057 ( .A(n981), .B(n976), .Y(n775) );
  CLKINVXL U1058 ( .A(n973), .Y(n875) );
  OAI22XL U1059 ( .A0(n36), .A1(n733), .B0(n732), .B1(n34), .Y(n598) );
  OAI22XL U1060 ( .A0(n12), .A1(n874), .B0(n9), .B1(n810), .Y(n562) );
  OAI22XL U1061 ( .A0(n42), .A1(n719), .B0(n718), .B1(n40), .Y(n584) );
  OAI22XL U1062 ( .A0(n42), .A1(n717), .B0(n716), .B1(n40), .Y(n582) );
  XNOR2XL U1063 ( .A(n981), .B(n977), .Y(n758) );
  OAI22XL U1064 ( .A0(n24), .A1(n761), .B0(n760), .B1(n22), .Y(n626) );
  XNOR2XL U1065 ( .A(n981), .B(n978), .Y(n741) );
  OAI22XL U1066 ( .A0(n36), .A1(n730), .B0(n729), .B1(n34), .Y(n595) );
  CLKINVXL U1067 ( .A(n979), .Y(n869) );
  NAND2BXL U1068 ( .AN(n981), .B(n977), .Y(n759) );
  INVX1 U1069 ( .A(n368), .Y(n369) );
  OAI22XL U1070 ( .A0(n42), .A1(n714), .B0(n713), .B1(n40), .Y(n579) );
  NAND2BXL U1071 ( .AN(n982), .B(n976), .Y(n776) );
  NAND2BXL U1072 ( .AN(n982), .B(n978), .Y(n742) );
  CLKINVXL U1073 ( .A(n743), .Y(n551) );
  CLKINVXL U1074 ( .A(n976), .Y(n872) );
  CLKINVXL U1075 ( .A(n978), .Y(n870) );
  CLKINVXL U1076 ( .A(n977), .Y(n871) );
  NAND2BXL U1077 ( .AN(n982), .B(n975), .Y(n793) );
  OAI22XL U1078 ( .A0(n42), .A1(n712), .B0(n711), .B1(n40), .Y(n577) );
  NAND2X4 U1079 ( .A(n958), .B(n867), .Y(n6) );
  XNOR2X1 U1080 ( .A(n980), .B(b[13]), .Y(n694) );
  OAI21X1 U1081 ( .A0(n52), .A1(n157), .B0(n158), .Y(n156) );
  CLKINVXL U1082 ( .A(n216), .Y(n321) );
  NOR2X1 U1083 ( .A(n157), .B(n124), .Y(n122) );
  INVX2 U1084 ( .A(n157), .Y(n159) );
  INVX2 U1085 ( .A(n158), .Y(n160) );
  AOI21XL U1086 ( .A0(n214), .A1(n234), .B0(n215), .Y(n213) );
  CLKINVXL U1087 ( .A(n211), .Y(n320) );
  OAI21XL U1088 ( .A0(n254), .A1(n241), .B0(n242), .Y(n240) );
  CLKINVXL U1089 ( .A(n238), .Y(n324) );
  NOR2BXL U1090 ( .AN(n221), .B(n216), .Y(n214) );
  CLKINVXL U1091 ( .A(n232), .Y(n323) );
  OAI21XL U1092 ( .A0(n224), .A1(n216), .B0(n219), .Y(n215) );
  CLKINVXL U1093 ( .A(n222), .Y(n224) );
  NAND2XL U1094 ( .A(n122), .B(n98), .Y(n96) );
  CLKINVXL U1095 ( .A(n233), .Y(n231) );
  OAI21XL U1096 ( .A0(n52), .A1(n120), .B0(n121), .Y(n119) );
  CLKINVXL U1097 ( .A(n123), .Y(n121) );
  NAND2X1 U1098 ( .A(n315), .B(n171), .Y(n61) );
  CLKINVXL U1099 ( .A(n53), .Y(n177) );
  OAI21XL U1100 ( .A0(n52), .A1(n170), .B0(n171), .Y(n169) );
  NAND2X1 U1101 ( .A(n316), .B(n184), .Y(n62) );
  CLKINVXL U1102 ( .A(n183), .Y(n316) );
  INVX2 U1103 ( .A(n246), .Y(n244) );
  OAI21X1 U1104 ( .A0(n271), .A1(n275), .B0(n272), .Y(n270) );
  NOR2X1 U1105 ( .A(n271), .B(n274), .Y(n269) );
  INVX2 U1106 ( .A(n166), .Y(n164) );
  XOR2X1 U1107 ( .A(n276), .B(n76), .Y(product[8]) );
  NAND2X1 U1108 ( .A(n330), .B(n275), .Y(n76) );
  INVX2 U1109 ( .A(n274), .Y(n330) );
  NAND2XL U1110 ( .A(n946), .B(n261), .Y(n73) );
  INVX2 U1111 ( .A(n248), .Y(n326) );
  NAND2X1 U1112 ( .A(n465), .B(n476), .Y(n239) );
  INVX2 U1113 ( .A(n266), .Y(n264) );
  NAND2XL U1114 ( .A(n389), .B(n398), .Y(n200) );
  NAND2X1 U1115 ( .A(n423), .B(n436), .Y(n219) );
  NAND2XL U1116 ( .A(n411), .B(n422), .Y(n212) );
  XOR2X1 U1117 ( .A(n254), .B(n72), .Y(product[12]) );
  NAND2XL U1118 ( .A(n326), .B(n249), .Y(n72) );
  NAND2X1 U1119 ( .A(n329), .B(n272), .Y(n75) );
  CLKINVXL U1120 ( .A(n194), .Y(n196) );
  INVX2 U1121 ( .A(n149), .Y(n151) );
  OAI21XL U1122 ( .A0(n52), .A1(n96), .B0(n97), .Y(n95) );
  INVX2 U1123 ( .A(n101), .Y(n99) );
  NOR2X1 U1124 ( .A(n53), .B(n87), .Y(n85) );
  OAI21XL U1125 ( .A0(n52), .A1(n87), .B0(n88), .Y(n86) );
  NAND2XL U1126 ( .A(n122), .B(n89), .Y(n87) );
  INVX2 U1127 ( .A(n100), .Y(n98) );
  AOI21XL U1128 ( .A0(n160), .A1(n135), .B0(n136), .Y(n134) );
  OAI21XL U1129 ( .A0(n149), .A1(n137), .B0(n140), .Y(n136) );
  NAND2X1 U1130 ( .A(n969), .B(n116), .Y(n56) );
  XOR2X2 U1131 ( .A(n106), .B(n55), .Y(product[29]) );
  NAND2X1 U1132 ( .A(n970), .B(n105), .Y(n55) );
  OAI21XL U1133 ( .A0(n52), .A1(n109), .B0(n110), .Y(n108) );
  ADDFX2 U1134 ( .A(n469), .B(n478), .CI(n467), .CO(n464), .S(n465) );
  NAND2X1 U1135 ( .A(n965), .B(n968), .Y(n278) );
  INVX2 U1136 ( .A(n283), .Y(n281) );
  NOR2X1 U1137 ( .A(n517), .B(n524), .Y(n271) );
  OAI21XL U1138 ( .A0(n140), .A1(n128), .B0(n129), .Y(n127) );
  AND2X1 U1139 ( .A(n945), .B(n302), .Y(n962) );
  NAND2X2 U1140 ( .A(n388), .B(n379), .Y(n191) );
  OR2X4 U1141 ( .A(n509), .B(n516), .Y(n964) );
  AOI21X1 U1142 ( .A0(n295), .A1(n967), .B0(n292), .Y(n290) );
  INVX2 U1143 ( .A(n294), .Y(n292) );
  OAI21X1 U1144 ( .A0(n298), .A1(n296), .B0(n297), .Y(n295) );
  AOI21X1 U1145 ( .A0(n945), .A1(n303), .B0(n300), .Y(n298) );
  INVX2 U1146 ( .A(n91), .Y(n308) );
  OAI21X1 U1147 ( .A0(n101), .A1(n91), .B0(n92), .Y(n90) );
  INVX2 U1148 ( .A(n105), .Y(n103) );
  INVX2 U1149 ( .A(n116), .Y(n114) );
  NAND2X1 U1150 ( .A(n969), .B(n970), .Y(n100) );
  NOR2X1 U1151 ( .A(n100), .B(n91), .Y(n89) );
  ADDFX2 U1152 ( .A(n535), .B(n538), .CI(n533), .CO(n530), .S(n531) );
  OR2XL U1153 ( .A(n691), .B(n563), .Y(n966) );
  ADDFX2 U1154 ( .A(n475), .B(n484), .CI(n473), .CO(n468), .S(n469) );
  ADDFX2 U1155 ( .A(n529), .B(n532), .CI(n527), .CO(n524), .S(n525) );
  OR2X1 U1156 ( .A(n541), .B(n544), .Y(n967) );
  NAND2X1 U1157 ( .A(n537), .B(n540), .Y(n288) );
  NAND2XL U1158 ( .A(n690), .B(n675), .Y(n305) );
  NAND2X1 U1159 ( .A(n541), .B(n544), .Y(n294) );
  NAND2X1 U1160 ( .A(n547), .B(n674), .Y(n302) );
  OR2X1 U1161 ( .A(n537), .B(n540), .Y(n968) );
  NAND2X1 U1162 ( .A(n350), .B(n347), .Y(n140) );
  NAND2XL U1163 ( .A(n346), .B(n343), .Y(n129) );
  OR2X1 U1164 ( .A(n342), .B(n341), .Y(n969) );
  NAND2X1 U1165 ( .A(n342), .B(n341), .Y(n116) );
  OR2X1 U1166 ( .A(n340), .B(n339), .Y(n970) );
  INVX2 U1167 ( .A(n338), .Y(n339) );
  NAND2X1 U1168 ( .A(n340), .B(n339), .Y(n105) );
  NOR2X1 U1169 ( .A(n564), .B(n338), .Y(n91) );
  NAND2X1 U1170 ( .A(n564), .B(n338), .Y(n92) );
  ADDFHX1 U1171 ( .A(n408), .B(n597), .CI(n642), .CO(n396), .S(n397) );
  OAI2BB1X1 U1172 ( .A0N(n16), .A1N(n18), .B0(n553), .Y(n642) );
  CLKINVXL U1173 ( .A(n777), .Y(n553) );
  ADDFHX1 U1174 ( .A(n386), .B(n580), .CI(n625), .CO(n376), .S(n377) );
  OAI2BB1X1 U1175 ( .A0N(n22), .A1N(n24), .B0(n552), .Y(n625) );
  INVX2 U1176 ( .A(n760), .Y(n552) );
  OAI2BB1X1 U1177 ( .A0N(n867), .A1N(n6), .B0(n555), .Y(n676) );
  OAI2BB1X1 U1178 ( .A0N(n9), .A1N(n12), .B0(n554), .Y(n659) );
  CLKINVXL U1179 ( .A(n794), .Y(n554) );
  ADDFHX1 U1180 ( .A(n583), .B(n598), .CI(n628), .CO(n404), .S(n405) );
  ADDFHX1 U1181 ( .A(n560), .B(n640), .CI(n670), .CO(n532), .S(n533) );
  OAI22XL U1182 ( .A0(n24), .A1(n775), .B0(n774), .B1(n22), .Y(n640) );
  INVX2 U1183 ( .A(n983), .Y(n981) );
  ADDFHX1 U1184 ( .A(n650), .B(n506), .CI(n497), .CO(n492), .S(n493) );
  NOR2BXL U1185 ( .AN(n981), .B(n40), .Y(n590) );
  INVX2 U1186 ( .A(n974), .Y(n874) );
  NOR2BXL U1187 ( .AN(n981), .B(n46), .Y(n573) );
  ADDFHX1 U1188 ( .A(n559), .B(n623), .CI(n638), .CO(n520), .S(n521) );
  CLKINVXL U1189 ( .A(n386), .Y(n387) );
  NOR2BXL U1190 ( .AN(n981), .B(n16), .Y(n658) );
  ADDHXL U1191 ( .A(n685), .B(n655), .CO(n534), .S(n535) );
  ADDFX2 U1192 ( .A(n354), .B(n576), .CI(n591), .CO(n348), .S(n349) );
  OAI2BB1X1 U1193 ( .A0N(n34), .A1N(n36), .B0(n550), .Y(n591) );
  INVX2 U1194 ( .A(n726), .Y(n550) );
  XNOR2X1 U1195 ( .A(n981), .B(n980), .Y(n707) );
  ADDHXL U1196 ( .A(n687), .B(n657), .CO(n542), .S(n543) );
  XNOR2X1 U1197 ( .A(n981), .B(n975), .Y(n792) );
  NOR2BXL U1198 ( .AN(n981), .B(n34), .Y(n607) );
  CMPR32X1 U1199 ( .A(n624), .B(n684), .C(n639), .CO(n528), .S(n529) );
  NOR2BXL U1200 ( .AN(n981), .B(n28), .Y(n624) );
  NOR2BXL U1201 ( .AN(n981), .B(n22), .Y(n641) );
  NAND2BX1 U1202 ( .AN(n982), .B(n980), .Y(n708) );
  INVX2 U1203 ( .A(n983), .Y(n982) );
  ADDFX2 U1204 ( .A(n575), .B(n345), .CI(n348), .CO(n342), .S(n343) );
  INVX2 U1205 ( .A(n344), .Y(n345) );
  OAI2BB1X1 U1206 ( .A0N(n28), .A1N(n30), .B0(n551), .Y(n608) );
  NOR2BXL U1207 ( .AN(n981), .B(n9), .Y(n675) );
  XNOR2X1 U1208 ( .A(n981), .B(n974), .Y(n809) );
  CLKINVXL U1209 ( .A(n354), .Y(n355) );
  NAND2BX1 U1210 ( .AN(n982), .B(n974), .Y(n810) );
  CLKINVXL U1211 ( .A(n811), .Y(n555) );
  INVX2 U1212 ( .A(n980), .Y(n868) );
  NOR2BXL U1213 ( .AN(n981), .B(n867), .Y(product[0]) );
  ADDFX2 U1214 ( .A(n344), .B(n565), .CI(n574), .CO(n340), .S(n341) );
  OAI2BB1X1 U1215 ( .A0N(n40), .A1N(n42), .B0(n549), .Y(n574) );
  INVX2 U1216 ( .A(n709), .Y(n549) );
  OAI2BB1X1 U1217 ( .A0N(n46), .A1N(n48), .B0(n548), .Y(n564) );
  INVX2 U1218 ( .A(n692), .Y(n548) );
  XOR2X1 U1219 ( .A(n980), .B(a[14]), .Y(n844) );
  XOR2X1 U1220 ( .A(n976), .B(a[6]), .Y(n848) );
  BUFX20 U1221 ( .A(a[5]), .Y(n975) );
  XOR2X1 U1222 ( .A(n977), .B(a[8]), .Y(n847) );
  XOR2X1 U1223 ( .A(n978), .B(a[10]), .Y(n846) );
  XOR2X1 U1224 ( .A(n975), .B(a[4]), .Y(n849) );
  XOR2X1 U1225 ( .A(n974), .B(a[2]), .Y(n850) );
  BUFX12 U1226 ( .A(a[1]), .Y(n973) );
  XNOR2X1 U1227 ( .A(n973), .B(b[9]), .Y(n817) );
  XNOR2X1 U1228 ( .A(n980), .B(b[7]), .Y(n700) );
  XNOR2X1 U1229 ( .A(n980), .B(b[1]), .Y(n706) );
  XNOR2X1 U1230 ( .A(n980), .B(b[4]), .Y(n703) );
  XNOR2X1 U1231 ( .A(n980), .B(b[3]), .Y(n704) );
  XNOR2X1 U1232 ( .A(n980), .B(b[2]), .Y(n705) );
  XNOR2X1 U1233 ( .A(n977), .B(b[8]), .Y(n750) );
  XNOR2X1 U1234 ( .A(n977), .B(b[7]), .Y(n751) );
  XNOR2X1 U1235 ( .A(n976), .B(b[10]), .Y(n765) );
  XNOR2X1 U1236 ( .A(n974), .B(b[14]), .Y(n795) );
  XNOR2X1 U1237 ( .A(n978), .B(b[8]), .Y(n733) );
  XNOR2X1 U1238 ( .A(n976), .B(b[9]), .Y(n766) );
  XNOR2X1 U1239 ( .A(n974), .B(b[12]), .Y(n797) );
  XNOR2X1 U1240 ( .A(n977), .B(b[6]), .Y(n752) );
  XNOR2X1 U1241 ( .A(n975), .B(b[9]), .Y(n783) );
  XNOR2X1 U1242 ( .A(n975), .B(b[12]), .Y(n780) );
  XNOR2X1 U1243 ( .A(n977), .B(b[9]), .Y(n749) );
  XNOR2X1 U1244 ( .A(n974), .B(b[13]), .Y(n796) );
  XNOR2X1 U1245 ( .A(n974), .B(b[11]), .Y(n798) );
  XNOR2X1 U1246 ( .A(n977), .B(b[11]), .Y(n747) );
  XNOR2X1 U1247 ( .A(n978), .B(b[7]), .Y(n734) );
  XNOR2X1 U1248 ( .A(n975), .B(b[11]), .Y(n781) );
  XNOR2X1 U1249 ( .A(n977), .B(b[5]), .Y(n753) );
  XNOR2X1 U1250 ( .A(n978), .B(b[9]), .Y(n732) );
  XNOR2X1 U1251 ( .A(n975), .B(b[13]), .Y(n779) );
  XNOR2X1 U1252 ( .A(n975), .B(b[14]), .Y(n778) );
  XNOR2X1 U1253 ( .A(n975), .B(b[8]), .Y(n784) );
  XNOR2X1 U1254 ( .A(n974), .B(b[10]), .Y(n799) );
  XNOR2X1 U1255 ( .A(n977), .B(b[10]), .Y(n748) );
  XNOR2X1 U1256 ( .A(n976), .B(b[6]), .Y(n769) );
  XNOR2X1 U1257 ( .A(n978), .B(b[1]), .Y(n740) );
  XNOR2X1 U1258 ( .A(n975), .B(b[5]), .Y(n787) );
  XNOR2X1 U1259 ( .A(n975), .B(b[6]), .Y(n786) );
  XNOR2X1 U1260 ( .A(n974), .B(b[9]), .Y(n800) );
  XNOR2X1 U1261 ( .A(n976), .B(b[4]), .Y(n771) );
  XNOR2X1 U1262 ( .A(n975), .B(b[7]), .Y(n785) );
  XNOR2X1 U1263 ( .A(n978), .B(b[4]), .Y(n737) );
  XNOR2X1 U1264 ( .A(n975), .B(b[10]), .Y(n782) );
  XNOR2X1 U1265 ( .A(n978), .B(b[2]), .Y(n739) );
  XNOR2X1 U1266 ( .A(n976), .B(b[5]), .Y(n770) );
  XNOR2X1 U1267 ( .A(n976), .B(b[8]), .Y(n767) );
  XNOR2X1 U1268 ( .A(n975), .B(b[4]), .Y(n788) );
  XNOR2X1 U1269 ( .A(n978), .B(b[10]), .Y(n731) );
  XNOR2X1 U1270 ( .A(n977), .B(b[3]), .Y(n755) );
  XNOR2X1 U1271 ( .A(n976), .B(b[7]), .Y(n768) );
  XNOR2X1 U1272 ( .A(n977), .B(b[1]), .Y(n757) );
  XNOR2X1 U1273 ( .A(n976), .B(b[3]), .Y(n772) );
  XNOR2X1 U1274 ( .A(n978), .B(b[3]), .Y(n738) );
  XNOR2X1 U1275 ( .A(n974), .B(b[3]), .Y(n806) );
  XNOR2X1 U1276 ( .A(n978), .B(b[12]), .Y(n729) );
  XNOR2X1 U1277 ( .A(n977), .B(b[4]), .Y(n754) );
  XNOR2X1 U1278 ( .A(n974), .B(b[2]), .Y(n807) );
  XNOR2X1 U1279 ( .A(n975), .B(b[3]), .Y(n789) );
  XNOR2X1 U1280 ( .A(n977), .B(b[2]), .Y(n756) );
  XNOR2X1 U1281 ( .A(n978), .B(b[11]), .Y(n730) );
  XNOR2X1 U1282 ( .A(n976), .B(b[1]), .Y(n774) );
  XNOR2X1 U1283 ( .A(n975), .B(b[1]), .Y(n791) );
  XNOR2X1 U1284 ( .A(n974), .B(b[1]), .Y(n808) );
  XNOR2X1 U1285 ( .A(n976), .B(b[14]), .Y(n761) );
  XNOR2X1 U1286 ( .A(n975), .B(b[2]), .Y(n790) );
  XNOR2X1 U1287 ( .A(n974), .B(b[6]), .Y(n803) );
  XNOR2X1 U1288 ( .A(n980), .B(b[9]), .Y(n698) );
  XNOR2X1 U1289 ( .A(n980), .B(b[8]), .Y(n699) );
  XNOR2X1 U1290 ( .A(n978), .B(b[5]), .Y(n736) );
  XNOR2X1 U1291 ( .A(n976), .B(b[2]), .Y(n773) );
  XNOR2X1 U1292 ( .A(n974), .B(b[5]), .Y(n804) );
  XNOR2X1 U1293 ( .A(n974), .B(b[8]), .Y(n801) );
  XNOR2X1 U1294 ( .A(n978), .B(b[6]), .Y(n735) );
  XNOR2X1 U1295 ( .A(n976), .B(b[12]), .Y(n763) );
  XNOR2X1 U1296 ( .A(n974), .B(b[4]), .Y(n805) );
  XNOR2X1 U1297 ( .A(n976), .B(b[11]), .Y(n764) );
  XNOR2X1 U1298 ( .A(n974), .B(b[7]), .Y(n802) );
  XNOR2X1 U1299 ( .A(n978), .B(b[13]), .Y(n728) );
  XNOR2X1 U1300 ( .A(n976), .B(b[13]), .Y(n762) );
  XNOR2X1 U1301 ( .A(n977), .B(b[14]), .Y(n744) );
  XNOR2X1 U1302 ( .A(n977), .B(b[12]), .Y(n746) );
  XNOR2X1 U1303 ( .A(n977), .B(b[13]), .Y(n745) );
  XNOR2X1 U1304 ( .A(n978), .B(b[14]), .Y(n727) );
  XNOR2XL U1305 ( .A(n980), .B(b[12]), .Y(n695) );
  XNOR2X1 U1306 ( .A(n980), .B(b[14]), .Y(n693) );
  OAI21X1 U1307 ( .A0(n254), .A1(n248), .B0(n249), .Y(n247) );
  OAI22XL U1308 ( .A0(n42), .A1(n722), .B0(n721), .B1(n40), .Y(n587) );
  CLKINVX4 U1309 ( .A(n51), .Y(n971) );
  INVX8 U1310 ( .A(n971), .Y(n972) );
  AOI21XL U1311 ( .A0(n972), .A1(n118), .B0(n119), .Y(n117) );
  XOR2X2 U1312 ( .A(n117), .B(n56), .Y(product[28]) );
  ADDFHX1 U1313 ( .A(n558), .B(n606), .CI(n666), .CO(n504), .S(n505) );
  XNOR2XL U1314 ( .A(n980), .B(b[15]), .Y(n692) );
  XNOR2X1 U1315 ( .A(n977), .B(b[15]), .Y(n743) );
  XNOR2X1 U1316 ( .A(n978), .B(b[15]), .Y(n726) );
  XNOR2X1 U1317 ( .A(n976), .B(b[15]), .Y(n760) );
  XNOR2X1 U1318 ( .A(n975), .B(b[15]), .Y(n777) );
  XNOR2X1 U1319 ( .A(n974), .B(b[15]), .Y(n794) );
  NOR2X4 U1320 ( .A(n437), .B(n450), .Y(n227) );
  ADDFHX2 U1321 ( .A(n636), .B(n621), .CI(n507), .CO(n502), .S(n503) );
  INVX2 U1322 ( .A(n268), .Y(n267) );
  OAI21X1 U1323 ( .A0(n304), .A1(n307), .B0(n305), .Y(n303) );
  XOR2XL U1324 ( .A(n82), .B(n307), .Y(product[2]) );
  NAND2XL U1325 ( .A(n691), .B(n563), .Y(n307) );
  XNOR2X1 U1326 ( .A(n973), .B(b[3]), .Y(n823) );
  NAND2BXL U1327 ( .AN(n981), .B(n973), .Y(n827) );
  XNOR2X1 U1328 ( .A(n973), .B(b[12]), .Y(n814) );
  XNOR2X1 U1329 ( .A(n973), .B(b[14]), .Y(n812) );
  XNOR2XL U1330 ( .A(n981), .B(n973), .Y(n826) );
  XNOR2X1 U1331 ( .A(n973), .B(b[13]), .Y(n813) );
  XNOR2X1 U1332 ( .A(n973), .B(b[4]), .Y(n822) );
  XNOR2X1 U1333 ( .A(n973), .B(b[5]), .Y(n821) );
  XNOR2X1 U1334 ( .A(n973), .B(b[15]), .Y(n811) );
  XNOR2X1 U1335 ( .A(n973), .B(b[10]), .Y(n816) );
  XNOR2X1 U1336 ( .A(n973), .B(b[6]), .Y(n820) );
  XNOR2X1 U1337 ( .A(n973), .B(b[8]), .Y(n818) );
  XNOR2X1 U1338 ( .A(n973), .B(b[11]), .Y(n815) );
  XNOR2X1 U1339 ( .A(n973), .B(b[7]), .Y(n819) );
  XNOR2X1 U1340 ( .A(n973), .B(b[1]), .Y(n825) );
  XNOR2X1 U1341 ( .A(n973), .B(b[2]), .Y(n824) );
  XNOR2X1 U1342 ( .A(n979), .B(b[15]), .Y(n709) );
  XNOR2X1 U1343 ( .A(n979), .B(b[14]), .Y(n710) );
  XNOR2X1 U1344 ( .A(n979), .B(b[13]), .Y(n711) );
  XNOR2X1 U1345 ( .A(n979), .B(b[12]), .Y(n712) );
  XNOR2X1 U1346 ( .A(n979), .B(b[11]), .Y(n713) );
  XNOR2X1 U1347 ( .A(n979), .B(b[9]), .Y(n715) );
  XNOR2X1 U1348 ( .A(n979), .B(b[10]), .Y(n714) );
  XNOR2X1 U1349 ( .A(n979), .B(b[8]), .Y(n716) );
  XNOR2X1 U1350 ( .A(n979), .B(b[7]), .Y(n717) );
  XNOR2X1 U1351 ( .A(n979), .B(b[6]), .Y(n718) );
  NAND2BXL U1352 ( .AN(n982), .B(n979), .Y(n725) );
  XNOR2X1 U1353 ( .A(n979), .B(b[5]), .Y(n719) );
  XNOR2XL U1354 ( .A(n981), .B(n979), .Y(n724) );
  XNOR2X1 U1355 ( .A(n979), .B(b[1]), .Y(n723) );
  XNOR2X1 U1356 ( .A(n979), .B(b[2]), .Y(n722) );
  XNOR2X1 U1357 ( .A(n979), .B(b[4]), .Y(n720) );
  XNOR2X1 U1358 ( .A(n979), .B(b[3]), .Y(n721) );
  XOR2X1 U1359 ( .A(n979), .B(a[12]), .Y(n845) );
  OAI21XL U1360 ( .A0(n196), .A1(n188), .B0(n191), .Y(n187) );
  INVX2 U1361 ( .A(n290), .Y(n289) );
  NAND2X1 U1362 ( .A(n209), .B(n221), .Y(n207) );
  XOR2X1 U1363 ( .A(n80), .B(n298), .Y(product[4]) );
endmodule


module PE_DW_mult_tc_29 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n6, n9, n12, n16, n18, n22, n24, n28, n30, n34, n36, n40, n42, n46,
         n48, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n62, n63, n64,
         n66, n67, n68, n70, n72, n73, n75, n76, n77, n79, n80, n82, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n103, n105, n106, n107, n108, n109, n110, n114, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n140, n141,
         n142, n143, n144, n145, n148, n149, n151, n154, n155, n156, n157,
         n158, n159, n160, n164, n166, n167, n168, n169, n170, n171, n173,
         n176, n177, n181, n182, n183, n184, n185, n186, n187, n188, n191,
         n192, n193, n194, n196, n199, n200, n201, n203, n204, n205, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n219, n220,
         n221, n222, n224, n227, n228, n229, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n244, n246, n247, n248,
         n249, n251, n254, n255, n256, n257, n259, n261, n262, n264, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n281, n283, n284, n286, n288, n289, n290, n292, n294,
         n295, n296, n297, n298, n300, n302, n303, n304, n305, n307, n308,
         n312, n313, n315, n316, n318, n319, n320, n321, n322, n323, n324,
         n326, n329, n330, n334, n336, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n844, n845, n846, n847, n848, n849, n850, n851, n867, n868, n869,
         n870, n871, n873, n874, n875, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993;

  AOI21X1 U60 ( .A0(n123), .A1(n89), .B0(n90), .Y(n88) );
  AOI21X1 U72 ( .A0(n123), .A1(n98), .B0(n99), .Y(n97) );
  AOI21X1 U76 ( .A0(n114), .A1(n983), .B0(n103), .Y(n101) );
  AOI21X1 U88 ( .A0(n123), .A1(n982), .B0(n114), .Y(n110) );
  AOI21X1 U106 ( .A0(n126), .A1(n151), .B0(n127), .Y(n125) );
  AOI21X1 U118 ( .A0(n160), .A1(n135), .B0(n136), .Y(n134) );
  AOI21X1 U132 ( .A0(n160), .A1(n313), .B0(n151), .Y(n145) );
  AOI21X1 U144 ( .A0(n51), .A1(n155), .B0(n156), .Y(n154) );
  AOI21X1 U194 ( .A0(n51), .A1(n193), .B0(n194), .Y(n192) );
  AOI21X1 U206 ( .A0(n51), .A1(n319), .B0(n203), .Y(n201) );
  AOI21X1 U216 ( .A0(n209), .A1(n222), .B0(n210), .Y(n208) );
  NOR2X2 U221 ( .A(n411), .B(n422), .Y(n211) );
  AOI21X1 U224 ( .A0(n214), .A1(n234), .B0(n215), .Y(n213) );
  NOR2X2 U231 ( .A(n423), .B(n436), .Y(n216) );
  AOI21X1 U234 ( .A0(n234), .A1(n221), .B0(n222), .Y(n220) );
  AOI21X1 U246 ( .A0(n234), .A1(n323), .B0(n231), .Y(n229) );
  NOR2X2 U251 ( .A(n451), .B(n464), .Y(n232) );
  NOR2X2 U256 ( .A(n241), .B(n238), .Y(n236) );
  AOI21X1 U294 ( .A0(n267), .A1(n976), .B0(n264), .Y(n262) );
  ADDFHX4 U385 ( .A(n382), .B(n373), .CI(n380), .CO(n370), .S(n371) );
  ADDFHX4 U408 ( .A(n629), .B(n614), .CI(n432), .CO(n416), .S(n417) );
  ADDFHX4 U411 ( .A(n427), .B(n438), .CI(n425), .CO(n422), .S(n423) );
  ADDFHX4 U418 ( .A(n441), .B(n452), .CI(n439), .CO(n436), .S(n437) );
  ADDFHX4 U419 ( .A(n456), .B(n443), .CI(n454), .CO(n438), .S(n439) );
  ADDFHX4 U421 ( .A(n462), .B(n449), .CI(n460), .CO(n442), .S(n443) );
  ADDFHX4 U426 ( .A(n455), .B(n466), .CI(n453), .CO(n450), .S(n451) );
  ADDFHX4 U427 ( .A(n461), .B(n457), .CI(n468), .CO(n452), .S(n453) );
  ADDFHX4 U445 ( .A(n493), .B(n500), .CI(n491), .CO(n488), .S(n489) );
  ADDFHX4 U450 ( .A(n503), .B(n510), .CI(n501), .CO(n498), .S(n499) );
  ADDFHX4 U451 ( .A(n514), .B(n512), .CI(n505), .CO(n500), .S(n501) );
  OAI22X1 U478 ( .A0(n48), .A1(n693), .B0(n46), .B1(n692), .Y(n338) );
  OAI22X1 U479 ( .A0(n48), .A1(n694), .B0(n46), .B1(n693), .Y(n565) );
  OAI22X1 U480 ( .A0(n48), .A1(n695), .B0(n46), .B1(n694), .Y(n344) );
  OAI22X1 U481 ( .A0(n48), .A1(n696), .B0(n46), .B1(n695), .Y(n566) );
  OAI22X1 U482 ( .A0(n48), .A1(n697), .B0(n46), .B1(n696), .Y(n354) );
  OAI22X1 U483 ( .A0(n48), .A1(n698), .B0(n46), .B1(n697), .Y(n567) );
  OAI22X1 U484 ( .A0(n48), .A1(n699), .B0(n46), .B1(n698), .Y(n368) );
  OAI22X1 U485 ( .A0(n48), .A1(n700), .B0(n46), .B1(n699), .Y(n568) );
  OAI22X1 U487 ( .A0(n48), .A1(n702), .B0(n46), .B1(n701), .Y(n569) );
  OAI22X1 U489 ( .A0(n48), .A1(n704), .B0(n46), .B1(n703), .Y(n570) );
  OAI22X1 U491 ( .A0(n48), .A1(n706), .B0(n46), .B1(n705), .Y(n571) );
  OAI22X1 U492 ( .A0(n48), .A1(n707), .B0(n46), .B1(n706), .Y(n572) );
  OAI22X1 U511 ( .A0(n42), .A1(n869), .B0(n40), .B1(n725), .Y(n557) );
  OAI22X1 U514 ( .A0(n42), .A1(n710), .B0(n709), .B1(n40), .Y(n575) );
  OAI22X1 U515 ( .A0(n42), .A1(n711), .B0(n710), .B1(n40), .Y(n576) );
  OAI22X1 U517 ( .A0(n42), .A1(n713), .B0(n712), .B1(n40), .Y(n578) );
  OAI22X1 U519 ( .A0(n42), .A1(n715), .B0(n714), .B1(n40), .Y(n580) );
  OAI22X1 U520 ( .A0(n42), .A1(n716), .B0(n715), .B1(n40), .Y(n581) );
  OAI22X1 U522 ( .A0(n42), .A1(n718), .B0(n717), .B1(n40), .Y(n583) );
  OAI22X1 U526 ( .A0(n42), .A1(n722), .B0(n721), .B1(n40), .Y(n587) );
  OAI22X1 U527 ( .A0(n42), .A1(n723), .B0(n722), .B1(n40), .Y(n588) );
  OAI22X1 U547 ( .A0(n36), .A1(n870), .B0(n34), .B1(n742), .Y(n558) );
  OAI22X1 U550 ( .A0(n36), .A1(n727), .B0(n726), .B1(n34), .Y(n592) );
  OAI22X1 U551 ( .A0(n36), .A1(n728), .B0(n727), .B1(n34), .Y(n593) );
  OAI22X1 U552 ( .A0(n36), .A1(n729), .B0(n728), .B1(n34), .Y(n594) );
  OAI22X1 U554 ( .A0(n36), .A1(n731), .B0(n730), .B1(n34), .Y(n596) );
  OAI22X1 U557 ( .A0(n36), .A1(n734), .B0(n733), .B1(n34), .Y(n599) );
  OAI22X1 U558 ( .A0(n36), .A1(n735), .B0(n734), .B1(n34), .Y(n600) );
  OAI22X1 U559 ( .A0(n36), .A1(n736), .B0(n735), .B1(n34), .Y(n601) );
  OAI22X1 U560 ( .A0(n36), .A1(n737), .B0(n736), .B1(n34), .Y(n602) );
  OAI22X1 U561 ( .A0(n36), .A1(n738), .B0(n737), .B1(n34), .Y(n603) );
  OAI22X1 U562 ( .A0(n36), .A1(n739), .B0(n738), .B1(n34), .Y(n604) );
  OAI22X1 U563 ( .A0(n36), .A1(n740), .B0(n739), .B1(n34), .Y(n605) );
  OAI22X1 U564 ( .A0(n36), .A1(n741), .B0(n740), .B1(n34), .Y(n606) );
  OAI22X1 U662 ( .A0(n18), .A1(n782), .B0(n781), .B1(n951), .Y(n647) );
  OAI22X1 U666 ( .A0(n18), .A1(n786), .B0(n785), .B1(n951), .Y(n651) );
  OAI22X1 U667 ( .A0(n18), .A1(n787), .B0(n786), .B1(n951), .Y(n652) );
  OAI22X1 U694 ( .A0(n12), .A1(n795), .B0(n794), .B1(n9), .Y(n660) );
  OAI22X1 U695 ( .A0(n12), .A1(n796), .B0(n795), .B1(n9), .Y(n661) );
  OAI22X1 U696 ( .A0(n12), .A1(n797), .B0(n796), .B1(n9), .Y(n662) );
  OAI22X1 U700 ( .A0(n12), .A1(n801), .B0(n800), .B1(n9), .Y(n666) );
  OAI22X1 U701 ( .A0(n12), .A1(n802), .B0(n801), .B1(n9), .Y(n667) );
  OAI22X1 U702 ( .A0(n12), .A1(n803), .B0(n802), .B1(n9), .Y(n668) );
  OAI22X1 U703 ( .A0(n12), .A1(n804), .B0(n803), .B1(n9), .Y(n669) );
  OAI22X1 U704 ( .A0(n12), .A1(n805), .B0(n804), .B1(n9), .Y(n670) );
  OAI22X1 U705 ( .A0(n12), .A1(n806), .B0(n805), .B1(n9), .Y(n671) );
  OAI22X1 U708 ( .A0(n12), .A1(n809), .B0(n808), .B1(n9), .Y(n674) );
  OAI22X1 U733 ( .A0(n6), .A1(n815), .B0(n814), .B1(n867), .Y(n680) );
  OAI22X1 U735 ( .A0(n6), .A1(n817), .B0(n816), .B1(n867), .Y(n682) );
  OAI22X1 U736 ( .A0(n6), .A1(n818), .B0(n817), .B1(n867), .Y(n683) );
  OAI22X1 U738 ( .A0(n6), .A1(n820), .B0(n819), .B1(n867), .Y(n685) );
  OAI22X1 U740 ( .A0(n6), .A1(n822), .B0(n821), .B1(n867), .Y(n687) );
  OAI22X1 U741 ( .A0(n6), .A1(n823), .B0(n822), .B1(n867), .Y(n688) );
  OAI22X1 U742 ( .A0(n6), .A1(n824), .B0(n823), .B1(n867), .Y(n689) );
  NAND2X4 U786 ( .A(n46), .B(n844), .Y(n48) );
  XNOR2X4 U788 ( .A(n992), .B(a[14]), .Y(n46) );
  NAND2X4 U789 ( .A(n40), .B(n845), .Y(n42) );
  XNOR2X4 U791 ( .A(n991), .B(a[12]), .Y(n40) );
  NAND2X4 U792 ( .A(n34), .B(n846), .Y(n36) );
  XNOR2X4 U794 ( .A(n990), .B(a[10]), .Y(n34) );
  NAND2X4 U795 ( .A(n28), .B(n847), .Y(n30) );
  NAND2X4 U798 ( .A(n953), .B(n848), .Y(n24) );
  XNOR2X4 U800 ( .A(n988), .B(a[6]), .Y(n22) );
  NAND2X4 U801 ( .A(n950), .B(n849), .Y(n18) );
  XNOR2X4 U803 ( .A(n987), .B(a[4]), .Y(n16) );
  NAND2X4 U804 ( .A(n9), .B(n850), .Y(n12) );
  XNOR2X4 U806 ( .A(n986), .B(a[2]), .Y(n9) );
  NAND2X4 U807 ( .A(n851), .B(n867), .Y(n6) );
  INVX4 U812 ( .A(n949), .Y(n951) );
  NOR2BXL U813 ( .AN(n193), .B(n188), .Y(n186) );
  NAND2BX1 U814 ( .AN(n188), .B(n191), .Y(n63) );
  XNOR2XL U815 ( .A(n993), .B(b[15]), .Y(n692) );
  XNOR2XL U816 ( .A(n992), .B(b[15]), .Y(n709) );
  XNOR2XL U817 ( .A(n991), .B(b[15]), .Y(n726) );
  ADDFHX1 U818 ( .A(n504), .B(n502), .CI(n495), .CO(n490), .S(n491) );
  ADDFHX1 U819 ( .A(n636), .B(n621), .CI(n507), .CO(n502), .S(n503) );
  XOR2X2 U820 ( .A(n192), .B(n63), .Y(product[21]) );
  BUFX12 U821 ( .A(a[5]), .Y(n988) );
  NOR2BX2 U822 ( .AN(b[0]), .B(n954), .Y(n641) );
  INVX3 U823 ( .A(n952), .Y(n954) );
  OAI22X1 U824 ( .A0(n6), .A1(n819), .B0(n818), .B1(n867), .Y(n684) );
  NAND2X4 U825 ( .A(n943), .B(n944), .Y(n945) );
  NAND2X4 U826 ( .A(n945), .B(n208), .Y(n51) );
  CLKINVX2 U827 ( .A(n207), .Y(n943) );
  INVX3 U828 ( .A(n235), .Y(n944) );
  NAND2X1 U829 ( .A(n209), .B(n221), .Y(n207) );
  AOI21X1 U830 ( .A0(n51), .A1(n186), .B0(n187), .Y(n185) );
  NOR2XL U831 ( .A(n30), .B(n756), .Y(n946) );
  NOR2XL U832 ( .A(n755), .B(n28), .Y(n947) );
  OR2X2 U833 ( .A(n946), .B(n947), .Y(n621) );
  OR2X4 U834 ( .A(n278), .B(n290), .Y(n948) );
  NAND2X4 U835 ( .A(n948), .B(n279), .Y(n277) );
  NAND2X2 U836 ( .A(n981), .B(n978), .Y(n278) );
  AOI21X4 U837 ( .A0(n295), .A1(n979), .B0(n292), .Y(n290) );
  AOI21X2 U838 ( .A0(n981), .A1(n286), .B0(n281), .Y(n279) );
  CLKINVX2 U839 ( .A(n277), .Y(n276) );
  INVX4 U840 ( .A(n16), .Y(n949) );
  CLKINVX4 U841 ( .A(n949), .Y(n950) );
  INVX4 U842 ( .A(n22), .Y(n952) );
  CLKINVX4 U843 ( .A(n952), .Y(n953) );
  AOI21X4 U844 ( .A0(n974), .A1(n251), .B0(n244), .Y(n242) );
  ADDFHX1 U845 ( .A(n641), .B(n686), .CI(n656), .CO(n538), .S(n539) );
  BUFX12 U846 ( .A(a[3]), .Y(n987) );
  OAI22X1 U847 ( .A0(n18), .A1(n788), .B0(n787), .B1(n951), .Y(n653) );
  AOI21XL U848 ( .A0(n51), .A1(n85), .B0(n86), .Y(product[31]) );
  AOI21XL U849 ( .A0(n51), .A1(n94), .B0(n95), .Y(n93) );
  AOI21XL U850 ( .A0(n51), .A1(n107), .B0(n108), .Y(n106) );
  AOI21XL U851 ( .A0(n51), .A1(n118), .B0(n119), .Y(n117) );
  AOI21XL U852 ( .A0(n51), .A1(n131), .B0(n132), .Y(n130) );
  AOI21XL U853 ( .A0(n51), .A1(n168), .B0(n169), .Y(n167) );
  AOI21XL U854 ( .A0(n51), .A1(n142), .B0(n143), .Y(n141) );
  NOR2X2 U855 ( .A(n465), .B(n476), .Y(n238) );
  ADDFHX2 U856 ( .A(n469), .B(n478), .CI(n467), .CO(n464), .S(n465) );
  AOI21X1 U857 ( .A0(n51), .A1(n177), .B0(n972), .Y(n176) );
  OAI21X2 U858 ( .A0(n242), .A1(n238), .B0(n239), .Y(n237) );
  AOI21X1 U859 ( .A0(n957), .A1(n264), .B0(n259), .Y(n257) );
  OAI22X1 U860 ( .A0(n18), .A1(n778), .B0(n777), .B1(n951), .Y(n643) );
  XNOR2X2 U861 ( .A(n986), .B(b[5]), .Y(n821) );
  CMPR32X1 U862 ( .A(n408), .B(n597), .C(n642), .CO(n396), .S(n397) );
  INVX1 U863 ( .A(n408), .Y(n409) );
  OAI22X2 U864 ( .A0(n48), .A1(n703), .B0(n46), .B1(n702), .Y(n408) );
  ADDFHX1 U865 ( .A(n558), .B(n606), .CI(n666), .CO(n504), .S(n505) );
  INVX1 U866 ( .A(n643), .Y(n955) );
  CLKINVX2 U867 ( .A(n955), .Y(n956) );
  ADDHX1 U868 ( .A(n681), .B(n651), .CO(n506), .S(n507) );
  XNOR2X2 U869 ( .A(n986), .B(b[6]), .Y(n820) );
  XNOR2X2 U870 ( .A(n988), .B(b[6]), .Y(n786) );
  OAI22X2 U871 ( .A0(n24), .A1(n771), .B0(n770), .B1(n954), .Y(n636) );
  NOR2X2 U872 ( .A(n389), .B(n398), .Y(n199) );
  ADDFHX2 U873 ( .A(n402), .B(n400), .CI(n391), .CO(n388), .S(n389) );
  ADDFHX1 U874 ( .A(n403), .B(n412), .CI(n401), .CO(n398), .S(n399) );
  ADDFHX1 U875 ( .A(n613), .B(n956), .CI(n409), .CO(n406), .S(n407) );
  XOR2X2 U876 ( .A(n989), .B(a[6]), .Y(n848) );
  XOR2X2 U877 ( .A(n988), .B(a[4]), .Y(n849) );
  XNOR2X2 U878 ( .A(n986), .B(b[11]), .Y(n815) );
  XNOR2X2 U879 ( .A(n990), .B(b[11]), .Y(n747) );
  XOR2X4 U880 ( .A(n991), .B(a[10]), .Y(n846) );
  CMPR32X1 U881 ( .A(n568), .B(n595), .C(n610), .CO(n374), .S(n375) );
  NAND2XL U882 ( .A(n509), .B(n516), .Y(n266) );
  BUFX12 U883 ( .A(a[13]), .Y(n992) );
  BUFX8 U884 ( .A(a[15]), .Y(n993) );
  ADDFHX1 U885 ( .A(n367), .B(n365), .CI(n372), .CO(n362), .S(n363) );
  NAND2X1 U886 ( .A(n370), .B(n363), .Y(n171) );
  CMPR32X1 U887 ( .A(n386), .B(n580), .C(n625), .CO(n376), .S(n377) );
  NAND2X1 U888 ( .A(n989), .B(a[8]), .Y(n961) );
  CMPR32X1 U889 ( .A(n567), .B(n593), .C(n366), .CO(n358), .S(n359) );
  OR2X2 U890 ( .A(n477), .B(n488), .Y(n974) );
  ADDFX2 U891 ( .A(n566), .B(n352), .CI(n349), .CO(n346), .S(n347) );
  XOR2X1 U892 ( .A(n262), .B(n73), .Y(product[11]) );
  OAI21X2 U893 ( .A0(n268), .A1(n256), .B0(n257), .Y(n255) );
  NAND2X1 U894 ( .A(n957), .B(n976), .Y(n256) );
  NAND2X1 U895 ( .A(n451), .B(n464), .Y(n233) );
  INVX2 U896 ( .A(n53), .Y(n177) );
  XOR2X1 U897 ( .A(n141), .B(n58), .Y(product[26]) );
  XOR2X1 U898 ( .A(n167), .B(n60), .Y(product[24]) );
  XOR2X1 U899 ( .A(n154), .B(n59), .Y(product[25]) );
  OAI22X1 U900 ( .A0(n30), .A1(n757), .B0(n756), .B1(n28), .Y(n622) );
  OR2X1 U901 ( .A(n24), .B(n775), .Y(n963) );
  ADDFX2 U902 ( .A(n637), .B(n652), .CI(n667), .CO(n512), .S(n513) );
  ADDFX2 U903 ( .A(n635), .B(n665), .CI(n620), .CO(n494), .S(n495) );
  ADDFX2 U904 ( .A(n650), .B(n506), .CI(n497), .CO(n492), .S(n493) );
  ADDFX2 U905 ( .A(n557), .B(n984), .CI(n634), .CO(n484), .S(n485) );
  ADDFX2 U906 ( .A(n618), .B(n985), .CI(n648), .CO(n472), .S(n473) );
  BUFX2 U907 ( .A(n663), .Y(n985) );
  ADDFX2 U908 ( .A(n633), .B(n603), .CI(n486), .CO(n470), .S(n471) );
  ADDFX2 U909 ( .A(n596), .B(n626), .CI(n387), .CO(n384), .S(n385) );
  ADDHXL U910 ( .A(n689), .B(n562), .CO(n546), .S(n547) );
  ADDHXL U911 ( .A(n687), .B(n657), .CO(n542), .S(n543) );
  ADDFX2 U912 ( .A(n669), .B(n654), .CI(n534), .CO(n526), .S(n527) );
  ADDFX2 U913 ( .A(n668), .B(n523), .CI(n528), .CO(n518), .S(n519) );
  ADDFX2 U914 ( .A(n559), .B(n623), .CI(n638), .CO(n520), .S(n521) );
  ADDFX2 U915 ( .A(n513), .B(n518), .CI(n511), .CO(n508), .S(n509) );
  ADDFX2 U916 ( .A(n487), .B(n496), .CI(n494), .CO(n480), .S(n481) );
  ADDFX2 U917 ( .A(n434), .B(n599), .CI(n659), .CO(n420), .S(n421) );
  ADDFX2 U918 ( .A(n645), .B(n585), .CI(n630), .CO(n430), .S(n431) );
  ADDFX2 U919 ( .A(n615), .B(n660), .CI(n435), .CO(n432), .S(n433) );
  ADDFX2 U920 ( .A(n600), .B(n448), .CI(n446), .CO(n428), .S(n429) );
  XNOR2X1 U921 ( .A(n631), .B(n571), .Y(n449) );
  ADDFX2 U922 ( .A(n662), .B(n463), .CI(n474), .CO(n456), .S(n457) );
  ADDFHX1 U923 ( .A(n475), .B(n484), .CI(n473), .CO(n468), .S(n469) );
  ADDFX2 U924 ( .A(n485), .B(n483), .CI(n492), .CO(n478), .S(n479) );
  ADDFHX1 U925 ( .A(n472), .B(n470), .CI(n459), .CO(n454), .S(n455) );
  ADDFX2 U926 ( .A(n482), .B(n471), .CI(n480), .CO(n466), .S(n467) );
  ADDFX2 U927 ( .A(n418), .B(n416), .CI(n414), .CO(n400), .S(n401) );
  ADDFX2 U928 ( .A(n420), .B(n405), .CI(n407), .CO(n402), .S(n403) );
  ADDFX2 U929 ( .A(n627), .B(n406), .CI(n404), .CO(n392), .S(n393) );
  ADDFX2 U930 ( .A(n395), .B(n397), .CI(n393), .CO(n390), .S(n391) );
  ADDFX2 U931 ( .A(n611), .B(n581), .CI(n396), .CO(n382), .S(n383) );
  ADDFX2 U932 ( .A(n394), .B(n385), .CI(n383), .CO(n380), .S(n381) );
  ADDFX2 U933 ( .A(n594), .B(n579), .CI(n369), .CO(n366), .S(n367) );
  ADDFX2 U934 ( .A(n384), .B(n377), .CI(n375), .CO(n372), .S(n373) );
  ADDFX2 U935 ( .A(n609), .B(n376), .CI(n374), .CO(n364), .S(n365) );
  ADDFX2 U936 ( .A(n592), .B(n577), .CI(n355), .CO(n352), .S(n353) );
  OR2X1 U937 ( .A(n547), .B(n674), .Y(n980) );
  ADDFX2 U938 ( .A(n535), .B(n538), .CI(n533), .CO(n530), .S(n531) );
  NOR2X1 U939 ( .A(n489), .B(n498), .Y(n248) );
  INVX2 U940 ( .A(n266), .Y(n264) );
  CMPR32X1 U941 ( .A(n481), .B(n490), .C(n479), .CO(n476), .S(n477) );
  ADDFX2 U942 ( .A(n458), .B(n447), .CI(n445), .CO(n440), .S(n441) );
  ADDFX2 U943 ( .A(n428), .B(n417), .CI(n426), .CO(n412), .S(n413) );
  ADDFX2 U944 ( .A(n430), .B(n421), .CI(n419), .CO(n414), .S(n415) );
  ADDFHX1 U945 ( .A(n442), .B(n429), .CI(n440), .CO(n424), .S(n425) );
  NAND2X1 U946 ( .A(n399), .B(n410), .Y(n205) );
  ADDFX2 U947 ( .A(n392), .B(n390), .CI(n381), .CO(n378), .S(n379) );
  NAND2X1 U948 ( .A(n159), .B(n313), .Y(n144) );
  NOR2X1 U949 ( .A(n148), .B(n137), .Y(n135) );
  NOR2X1 U950 ( .A(n356), .B(n351), .Y(n148) );
  ADDFX2 U951 ( .A(n361), .B(n359), .CI(n364), .CO(n356), .S(n357) );
  ADDFX2 U952 ( .A(n360), .B(n353), .CI(n358), .CO(n350), .S(n351) );
  ADDFX2 U953 ( .A(n575), .B(n345), .CI(n348), .CO(n342), .S(n343) );
  NOR2X1 U954 ( .A(n690), .B(n675), .Y(n304) );
  XOR2X1 U955 ( .A(n267), .B(n968), .Y(product[10]) );
  XOR2X1 U956 ( .A(n993), .B(a[14]), .Y(n844) );
  NOR2X1 U957 ( .A(n137), .B(n128), .Y(n126) );
  AOI21X1 U958 ( .A0(n975), .A1(n173), .B0(n164), .Y(n158) );
  INVX2 U959 ( .A(n171), .Y(n173) );
  NOR2X1 U960 ( .A(n378), .B(n371), .Y(n183) );
  NOR2X1 U961 ( .A(n399), .B(n410), .Y(n204) );
  ADDFHX1 U962 ( .A(n415), .B(n424), .CI(n413), .CO(n410), .S(n411) );
  NOR2X1 U963 ( .A(n388), .B(n379), .Y(n188) );
  NAND2X1 U964 ( .A(n388), .B(n379), .Y(n191) );
  NOR2X1 U965 ( .A(n350), .B(n347), .Y(n137) );
  NOR2X1 U966 ( .A(n346), .B(n343), .Y(n128) );
  NOR2X1 U967 ( .A(n370), .B(n363), .Y(n170) );
  OR2X1 U968 ( .A(n362), .B(n357), .Y(n975) );
  NAND2X1 U969 ( .A(n356), .B(n351), .Y(n149) );
  XOR2X1 U970 ( .A(n284), .B(n77), .Y(product[7]) );
  NAND2X1 U971 ( .A(n321), .B(n219), .Y(n67) );
  XOR2X1 U972 ( .A(n229), .B(n68), .Y(product[16]) );
  NAND2X1 U973 ( .A(n122), .B(n982), .Y(n109) );
  OAI2BB1X1 U974 ( .A0N(n194), .A1N(n181), .B0(n973), .Y(n972) );
  INVX2 U975 ( .A(n182), .Y(n973) );
  OAI21X1 U976 ( .A0(n183), .A1(n191), .B0(n184), .Y(n182) );
  NOR2X1 U977 ( .A(n188), .B(n183), .Y(n181) );
  NAND2X1 U978 ( .A(n193), .B(n181), .Y(n53) );
  NOR2X1 U979 ( .A(n211), .B(n216), .Y(n209) );
  INVX2 U980 ( .A(a[0]), .Y(n867) );
  ADDFHX1 U981 ( .A(n607), .B(n682), .CI(n622), .CO(n514), .S(n515) );
  AOI21X2 U982 ( .A0(n269), .A1(n277), .B0(n270), .Y(n268) );
  OR2X4 U983 ( .A(n499), .B(n508), .Y(n957) );
  INVX2 U984 ( .A(n972), .Y(n52) );
  OR2X1 U985 ( .A(n691), .B(n563), .Y(n958) );
  BUFX8 U986 ( .A(a[7]), .Y(n989) );
  OAI22XL U987 ( .A0(n24), .A1(n762), .B0(n761), .B1(n954), .Y(n627) );
  OAI22XL U988 ( .A0(n24), .A1(n761), .B0(n760), .B1(n954), .Y(n626) );
  OAI22XL U989 ( .A0(n24), .A1(n763), .B0(n762), .B1(n954), .Y(n628) );
  OAI22XL U990 ( .A0(n24), .A1(n764), .B0(n763), .B1(n954), .Y(n629) );
  OAI22XL U991 ( .A0(n24), .A1(n765), .B0(n764), .B1(n954), .Y(n630) );
  OAI22XL U992 ( .A0(n24), .A1(n767), .B0(n766), .B1(n954), .Y(n632) );
  OAI22XL U993 ( .A0(n24), .A1(n769), .B0(n768), .B1(n954), .Y(n634) );
  OAI22XL U994 ( .A0(n24), .A1(n773), .B0(n772), .B1(n954), .Y(n638) );
  OAI22XL U995 ( .A0(n24), .A1(n770), .B0(n769), .B1(n954), .Y(n635) );
  OAI22XL U996 ( .A0(n24), .A1(n768), .B0(n767), .B1(n954), .Y(n633) );
  OAI22XL U997 ( .A0(n24), .A1(n774), .B0(n773), .B1(n954), .Y(n639) );
  OAI22XL U998 ( .A0(n24), .A1(n772), .B0(n771), .B1(n954), .Y(n637) );
  OAI22XL U999 ( .A0(n24), .A1(n766), .B0(n765), .B1(n954), .Y(n631) );
  NAND2X2 U1000 ( .A(n959), .B(n960), .Y(n962) );
  NAND2X4 U1001 ( .A(n961), .B(n962), .Y(n28) );
  INVX2 U1002 ( .A(n989), .Y(n959) );
  INVXL U1003 ( .A(a[8]), .Y(n960) );
  OAI22XL U1004 ( .A0(n30), .A1(n751), .B0(n750), .B1(n28), .Y(n616) );
  OAI22XL U1005 ( .A0(n30), .A1(n750), .B0(n749), .B1(n28), .Y(n615) );
  OAI22XL U1006 ( .A0(n30), .A1(n754), .B0(n753), .B1(n28), .Y(n619) );
  OAI22XL U1007 ( .A0(n30), .A1(n748), .B0(n747), .B1(n28), .Y(n613) );
  OAI22XL U1008 ( .A0(n30), .A1(n755), .B0(n754), .B1(n28), .Y(n620) );
  OAI22XL U1009 ( .A0(n30), .A1(n746), .B0(n745), .B1(n28), .Y(n611) );
  OAI22XL U1010 ( .A0(n30), .A1(n744), .B0(n743), .B1(n28), .Y(n609) );
  OAI22XL U1011 ( .A0(n30), .A1(n753), .B0(n752), .B1(n28), .Y(n618) );
  OAI22XL U1012 ( .A0(n30), .A1(n871), .B0(n28), .B1(n759), .Y(n559) );
  OAI22XL U1013 ( .A0(n30), .A1(n752), .B0(n751), .B1(n28), .Y(n617) );
  OAI22XL U1014 ( .A0(n30), .A1(n749), .B0(n748), .B1(n28), .Y(n614) );
  OAI22XL U1015 ( .A0(n30), .A1(n747), .B0(n746), .B1(n28), .Y(n612) );
  OAI22XL U1016 ( .A0(n30), .A1(n745), .B0(n744), .B1(n28), .Y(n610) );
  OR2X1 U1017 ( .A(n774), .B(n954), .Y(n964) );
  NAND2X2 U1018 ( .A(n963), .B(n964), .Y(n640) );
  XNOR2XL U1019 ( .A(b[0]), .B(n989), .Y(n775) );
  XNOR2X1 U1020 ( .A(n240), .B(n70), .Y(product[14]) );
  OAI21X1 U1021 ( .A0(n199), .A1(n205), .B0(n200), .Y(n194) );
  NOR2X1 U1022 ( .A(n204), .B(n199), .Y(n193) );
  INVX2 U1023 ( .A(n170), .Y(n315) );
  CLKINVXL U1024 ( .A(n238), .Y(n324) );
  INVX1 U1025 ( .A(n290), .Y(n289) );
  INVX2 U1026 ( .A(n148), .Y(n313) );
  OAI21X1 U1027 ( .A0(n158), .A1(n124), .B0(n125), .Y(n123) );
  INVX1 U1028 ( .A(n122), .Y(n120) );
  OAI21X2 U1029 ( .A0(n227), .A1(n233), .B0(n228), .Y(n222) );
  NOR2X1 U1030 ( .A(n227), .B(n232), .Y(n221) );
  NAND2X1 U1031 ( .A(n315), .B(n975), .Y(n157) );
  CLKINVX1 U1032 ( .A(n283), .Y(n281) );
  OR2X4 U1033 ( .A(n531), .B(n536), .Y(n981) );
  AOI21X1 U1034 ( .A0(n289), .A1(n978), .B0(n286), .Y(n284) );
  ADDFX2 U1035 ( .A(n354), .B(n576), .CI(n591), .CO(n348), .S(n349) );
  NAND2X1 U1036 ( .A(n437), .B(n450), .Y(n228) );
  NAND2X1 U1037 ( .A(n974), .B(n326), .Y(n241) );
  INVX1 U1038 ( .A(n248), .Y(n326) );
  INVX2 U1039 ( .A(n249), .Y(n251) );
  NAND2XL U1040 ( .A(n313), .B(n126), .Y(n124) );
  NAND2X1 U1041 ( .A(n159), .B(n135), .Y(n133) );
  NAND2X1 U1042 ( .A(n499), .B(n508), .Y(n261) );
  INVX1 U1043 ( .A(n288), .Y(n286) );
  XOR2X1 U1044 ( .A(n80), .B(n298), .Y(product[4]) );
  NAND2X1 U1045 ( .A(n334), .B(n297), .Y(n80) );
  OAI21X1 U1046 ( .A0(n140), .A1(n128), .B0(n129), .Y(n127) );
  NAND2XL U1047 ( .A(n981), .B(n283), .Y(n77) );
  XOR2XL U1048 ( .A(n82), .B(n307), .Y(product[2]) );
  ADDFHX2 U1049 ( .A(n521), .B(n526), .CI(n519), .CO(n516), .S(n517) );
  NAND2X1 U1050 ( .A(n690), .B(n675), .Y(n305) );
  ADDFHX1 U1051 ( .A(n670), .B(n640), .CI(n560), .CO(n532), .S(n533) );
  ADDFHX2 U1052 ( .A(n671), .B(n542), .CI(n539), .CO(n536), .S(n537) );
  INVX1 U1053 ( .A(n434), .Y(n435) );
  ADDFX2 U1054 ( .A(n619), .B(n589), .CI(n604), .CO(n482), .S(n483) );
  CLKINVXL U1055 ( .A(n386), .Y(n387) );
  INVX1 U1056 ( .A(n354), .Y(n355) );
  CLKINVXL U1057 ( .A(n811), .Y(n555) );
  BUFX20 U1058 ( .A(a[1]), .Y(n986) );
  BUFX20 U1059 ( .A(a[9]), .Y(n990) );
  BUFX20 U1060 ( .A(a[11]), .Y(n991) );
  INVX3 U1061 ( .A(n235), .Y(n234) );
  NAND2X1 U1062 ( .A(n324), .B(n239), .Y(n70) );
  XOR2X1 U1063 ( .A(n234), .B(n965), .Y(product[15]) );
  AND2X1 U1064 ( .A(n323), .B(n233), .Y(n965) );
  XOR2X1 U1065 ( .A(n220), .B(n67), .Y(product[17]) );
  XOR2X1 U1066 ( .A(n213), .B(n66), .Y(product[18]) );
  NAND2XL U1067 ( .A(n320), .B(n212), .Y(n66) );
  OAI21XL U1068 ( .A0(n52), .A1(n157), .B0(n158), .Y(n156) );
  OAI21XL U1069 ( .A0(n52), .A1(n144), .B0(n145), .Y(n143) );
  NOR2XL U1070 ( .A(n53), .B(n133), .Y(n131) );
  XOR2X1 U1071 ( .A(n185), .B(n62), .Y(product[22]) );
  NAND2XL U1072 ( .A(n316), .B(n184), .Y(n62) );
  XOR2X2 U1073 ( .A(n176), .B(n966), .Y(product[23]) );
  NAND2XL U1074 ( .A(n315), .B(n171), .Y(n966) );
  NAND2X2 U1075 ( .A(n423), .B(n436), .Y(n219) );
  XOR2X1 U1076 ( .A(n247), .B(n967), .Y(product[13]) );
  AND2X1 U1077 ( .A(n974), .B(n246), .Y(n967) );
  NAND2X1 U1078 ( .A(n465), .B(n476), .Y(n239) );
  XOR2X1 U1079 ( .A(n254), .B(n72), .Y(product[12]) );
  NAND2XL U1080 ( .A(n975), .B(n166), .Y(n60) );
  AND2X1 U1081 ( .A(n976), .B(n266), .Y(n968) );
  NAND2XL U1082 ( .A(n313), .B(n149), .Y(n59) );
  XNOR2X1 U1083 ( .A(n273), .B(n75), .Y(product[9]) );
  NAND2XL U1084 ( .A(n329), .B(n272), .Y(n75) );
  CLKINVXL U1085 ( .A(n271), .Y(n329) );
  NAND2XL U1086 ( .A(n389), .B(n398), .Y(n200) );
  NAND2XL U1087 ( .A(n330), .B(n275), .Y(n76) );
  CLKINVXL U1088 ( .A(n274), .Y(n330) );
  OR2X4 U1089 ( .A(n509), .B(n516), .Y(n976) );
  NAND2XL U1090 ( .A(n477), .B(n488), .Y(n246) );
  NAND2BX1 U1091 ( .AN(n128), .B(n129), .Y(n57) );
  XNOR2XL U1092 ( .A(n969), .B(n303), .Y(product[3]) );
  NAND2X1 U1093 ( .A(n980), .B(n302), .Y(n969) );
  XNOR2XL U1094 ( .A(n79), .B(n295), .Y(product[5]) );
  NAND2XL U1095 ( .A(n979), .B(n294), .Y(n79) );
  CLKINVXL U1096 ( .A(n296), .Y(n334) );
  CLKINVXL U1097 ( .A(n304), .Y(n336) );
  NAND2XL U1098 ( .A(n362), .B(n357), .Y(n166) );
  ADDFHX1 U1099 ( .A(n444), .B(n433), .CI(n431), .CO(n426), .S(n427) );
  ADDFX1 U1100 ( .A(n529), .B(n532), .CI(n527), .CO(n524), .S(n525) );
  NAND2XL U1101 ( .A(n531), .B(n536), .Y(n283) );
  NAND2X1 U1102 ( .A(n691), .B(n563), .Y(n307) );
  NAND2XL U1103 ( .A(n547), .B(n674), .Y(n302) );
  AND2X1 U1104 ( .A(n958), .B(n307), .Y(product[1]) );
  ADDFHX1 U1105 ( .A(n590), .B(n680), .CI(n605), .CO(n496), .S(n497) );
  OAI22XL U1106 ( .A0(n48), .A1(n868), .B0(n46), .B1(n708), .Y(n556) );
  OAI22XL U1107 ( .A0(n30), .A1(n758), .B0(n757), .B1(n28), .Y(n623) );
  OAI22XL U1108 ( .A0(n42), .A1(n721), .B0(n720), .B1(n40), .Y(n586) );
  OAI22XL U1109 ( .A0(n12), .A1(n800), .B0(n799), .B1(n9), .Y(n665) );
  OAI22XL U1110 ( .A0(n6), .A1(n816), .B0(n815), .B1(n867), .Y(n681) );
  OAI22XL U1111 ( .A0(n42), .A1(n724), .B0(n723), .B1(n40), .Y(n589) );
  CLKINVXL U1112 ( .A(n794), .Y(n554) );
  CLKINVXL U1113 ( .A(n777), .Y(n553) );
  OAI22XL U1114 ( .A0(n36), .A1(n732), .B0(n731), .B1(n34), .Y(n597) );
  ADDFX1 U1115 ( .A(n561), .B(n672), .CI(n543), .CO(n540), .S(n541) );
  CMPR32X1 U1116 ( .A(n658), .B(n688), .C(n673), .CO(n544), .S(n545) );
  OAI22XL U1117 ( .A0(n12), .A1(n808), .B0(n807), .B1(n9), .Y(n673) );
  OAI22XL U1118 ( .A0(n18), .A1(n792), .B0(n791), .B1(n951), .Y(n657) );
  OAI22XL U1119 ( .A0(n42), .A1(n720), .B0(n719), .B1(n40), .Y(n585) );
  OAI22XL U1120 ( .A0(n6), .A1(n812), .B0(n811), .B1(n867), .Y(n677) );
  OAI22XL U1121 ( .A0(n36), .A1(n733), .B0(n732), .B1(n34), .Y(n598) );
  XNOR2XL U1122 ( .A(b[0]), .B(n992), .Y(n724) );
  CLKINVXL U1123 ( .A(n760), .Y(n552) );
  OAI22XL U1124 ( .A0(n42), .A1(n719), .B0(n718), .B1(n40), .Y(n584) );
  NAND2BXL U1125 ( .AN(b[0]), .B(n989), .Y(n776) );
  OAI22XL U1126 ( .A0(n42), .A1(n717), .B0(n716), .B1(n40), .Y(n582) );
  NAND2BXL U1127 ( .AN(b[0]), .B(n992), .Y(n725) );
  NAND2BX1 U1128 ( .AN(b[0]), .B(n991), .Y(n742) );
  OAI22XL U1129 ( .A0(n36), .A1(n730), .B0(n729), .B1(n34), .Y(n595) );
  CLKINVXL U1130 ( .A(n992), .Y(n869) );
  NAND2BX1 U1131 ( .AN(b[0]), .B(n988), .Y(n793) );
  OAI22XL U1132 ( .A0(n42), .A1(n714), .B0(n713), .B1(n40), .Y(n579) );
  OAI22XL U1133 ( .A0(n42), .A1(n712), .B0(n711), .B1(n40), .Y(n577) );
  XNOR2X1 U1134 ( .A(n987), .B(b[14]), .Y(n795) );
  XNOR2X1 U1135 ( .A(n993), .B(b[3]), .Y(n704) );
  XNOR2X1 U1136 ( .A(n993), .B(b[1]), .Y(n706) );
  XNOR2X1 U1137 ( .A(n993), .B(b[2]), .Y(n705) );
  XNOR2X1 U1138 ( .A(n987), .B(b[11]), .Y(n798) );
  XNOR2X1 U1139 ( .A(n993), .B(b[5]), .Y(n702) );
  XNOR2X1 U1140 ( .A(n993), .B(b[7]), .Y(n700) );
  XNOR2X1 U1141 ( .A(n993), .B(b[4]), .Y(n703) );
  XNOR2X1 U1142 ( .A(n993), .B(b[6]), .Y(n701) );
  XNOR2X1 U1143 ( .A(n993), .B(b[8]), .Y(n699) );
  XNOR2X1 U1144 ( .A(n990), .B(b[14]), .Y(n744) );
  XNOR2X1 U1145 ( .A(n993), .B(b[9]), .Y(n698) );
  XNOR2X1 U1146 ( .A(n993), .B(b[11]), .Y(n696) );
  XNOR2X1 U1147 ( .A(n993), .B(b[10]), .Y(n697) );
  XNOR2X1 U1148 ( .A(n993), .B(b[13]), .Y(n694) );
  XNOR2X1 U1149 ( .A(n993), .B(b[12]), .Y(n695) );
  XNOR2X1 U1150 ( .A(n993), .B(b[14]), .Y(n693) );
  NOR2X1 U1151 ( .A(n53), .B(n144), .Y(n142) );
  NOR2X1 U1152 ( .A(n53), .B(n96), .Y(n94) );
  XOR2X2 U1153 ( .A(n201), .B(n64), .Y(product[20]) );
  NAND2X1 U1154 ( .A(n318), .B(n200), .Y(n64) );
  INVX2 U1155 ( .A(n199), .Y(n318) );
  CLKINVXL U1156 ( .A(n216), .Y(n321) );
  NAND2X1 U1157 ( .A(n322), .B(n228), .Y(n68) );
  CLKINVXL U1158 ( .A(n227), .Y(n322) );
  CLKINVXL U1159 ( .A(n211), .Y(n320) );
  INVX2 U1160 ( .A(n268), .Y(n267) );
  NOR2X1 U1161 ( .A(n157), .B(n124), .Y(n122) );
  OAI21X1 U1162 ( .A0(n254), .A1(n241), .B0(n242), .Y(n240) );
  INVX2 U1163 ( .A(n255), .Y(n254) );
  XOR2X1 U1164 ( .A(n51), .B(n971), .Y(product[19]) );
  AND2X1 U1165 ( .A(n319), .B(n205), .Y(n971) );
  INVX2 U1166 ( .A(n158), .Y(n160) );
  NOR2BXL U1167 ( .AN(n221), .B(n216), .Y(n214) );
  INVX2 U1168 ( .A(n157), .Y(n159) );
  CLKINVXL U1169 ( .A(n232), .Y(n323) );
  CLKINVXL U1170 ( .A(n222), .Y(n224) );
  CLKINVXL U1171 ( .A(n204), .Y(n319) );
  CLKINVXL U1172 ( .A(n233), .Y(n231) );
  CLKINVXL U1173 ( .A(n205), .Y(n203) );
  NAND2XL U1174 ( .A(n122), .B(n98), .Y(n96) );
  NOR2XL U1175 ( .A(n53), .B(n157), .Y(n155) );
  CLKINVXL U1176 ( .A(n183), .Y(n316) );
  INVX2 U1177 ( .A(n261), .Y(n259) );
  OAI21XL U1178 ( .A0(n52), .A1(n170), .B0(n171), .Y(n169) );
  NOR2XL U1179 ( .A(n53), .B(n170), .Y(n168) );
  INVX2 U1180 ( .A(n246), .Y(n244) );
  NAND2X1 U1181 ( .A(n411), .B(n422), .Y(n212) );
  XOR2X1 U1182 ( .A(n276), .B(n76), .Y(product[8]) );
  OAI21XL U1183 ( .A0(n52), .A1(n120), .B0(n121), .Y(n119) );
  INVX2 U1184 ( .A(n123), .Y(n121) );
  OAI21X1 U1185 ( .A0(n271), .A1(n275), .B0(n272), .Y(n270) );
  NOR2X1 U1186 ( .A(n271), .B(n274), .Y(n269) );
  NAND2X1 U1187 ( .A(n957), .B(n261), .Y(n73) );
  OAI21X1 U1188 ( .A0(n254), .A1(n248), .B0(n249), .Y(n247) );
  INVX2 U1189 ( .A(n166), .Y(n164) );
  NAND2XL U1190 ( .A(n326), .B(n249), .Y(n72) );
  INVX2 U1191 ( .A(n149), .Y(n151) );
  OAI21XL U1192 ( .A0(n276), .A1(n274), .B0(n275), .Y(n273) );
  OAI21XL U1193 ( .A0(n196), .A1(n188), .B0(n191), .Y(n187) );
  CLKINVXL U1194 ( .A(n194), .Y(n196) );
  OAI21XL U1195 ( .A0(n52), .A1(n96), .B0(n97), .Y(n95) );
  INVX2 U1196 ( .A(n101), .Y(n99) );
  NOR2X1 U1197 ( .A(n53), .B(n87), .Y(n85) );
  OAI21XL U1198 ( .A0(n52), .A1(n87), .B0(n88), .Y(n86) );
  NAND2XL U1199 ( .A(n122), .B(n89), .Y(n87) );
  INVX2 U1200 ( .A(n100), .Y(n98) );
  NAND2X1 U1201 ( .A(n312), .B(n140), .Y(n58) );
  CLKINVXL U1202 ( .A(n137), .Y(n312) );
  OAI21XL U1203 ( .A0(n52), .A1(n133), .B0(n134), .Y(n132) );
  OAI21XL U1204 ( .A0(n149), .A1(n137), .B0(n140), .Y(n136) );
  NAND2X1 U1205 ( .A(n983), .B(n105), .Y(n55) );
  NOR2XL U1206 ( .A(n53), .B(n109), .Y(n107) );
  OAI21XL U1207 ( .A0(n52), .A1(n109), .B0(n110), .Y(n108) );
  XOR2X2 U1208 ( .A(n117), .B(n56), .Y(product[28]) );
  NAND2X1 U1209 ( .A(n982), .B(n116), .Y(n56) );
  NOR2XL U1210 ( .A(n53), .B(n120), .Y(n118) );
  NOR2X1 U1211 ( .A(n525), .B(n530), .Y(n274) );
  NOR2X1 U1212 ( .A(n517), .B(n524), .Y(n271) );
  NAND2X2 U1213 ( .A(n489), .B(n498), .Y(n249) );
  INVX2 U1214 ( .A(n294), .Y(n292) );
  OAI21X1 U1215 ( .A0(n298), .A1(n296), .B0(n297), .Y(n295) );
  AOI21X1 U1216 ( .A0(n980), .A1(n303), .B0(n300), .Y(n298) );
  INVX2 U1217 ( .A(n302), .Y(n300) );
  NAND2X1 U1218 ( .A(n336), .B(n305), .Y(n82) );
  NAND2X1 U1219 ( .A(n517), .B(n524), .Y(n272) );
  XOR2X1 U1220 ( .A(n977), .B(n289), .Y(product[6]) );
  AND2X1 U1221 ( .A(n978), .B(n288), .Y(n977) );
  NAND2X1 U1222 ( .A(n378), .B(n371), .Y(n184) );
  OAI21X1 U1223 ( .A0(n304), .A1(n307), .B0(n305), .Y(n303) );
  NAND2X1 U1224 ( .A(n525), .B(n530), .Y(n275) );
  XOR2X1 U1225 ( .A(n93), .B(n54), .Y(product[30]) );
  NAND2X1 U1226 ( .A(n308), .B(n92), .Y(n54) );
  INVX2 U1227 ( .A(n91), .Y(n308) );
  OAI21X1 U1228 ( .A0(n101), .A1(n91), .B0(n92), .Y(n90) );
  INVX2 U1229 ( .A(n105), .Y(n103) );
  INVX2 U1230 ( .A(n116), .Y(n114) );
  NAND2X1 U1231 ( .A(n982), .B(n983), .Y(n100) );
  NOR2X1 U1232 ( .A(n100), .B(n91), .Y(n89) );
  ADDFX2 U1233 ( .A(n522), .B(n515), .CI(n520), .CO(n510), .S(n511) );
  OR2X1 U1234 ( .A(n537), .B(n540), .Y(n978) );
  OR2X1 U1235 ( .A(n541), .B(n544), .Y(n979) );
  NOR2X1 U1236 ( .A(n545), .B(n546), .Y(n296) );
  NAND2X1 U1237 ( .A(n537), .B(n540), .Y(n288) );
  NAND2X1 U1238 ( .A(n541), .B(n544), .Y(n294) );
  NAND2X1 U1239 ( .A(n545), .B(n546), .Y(n297) );
  NAND2X1 U1240 ( .A(n350), .B(n347), .Y(n140) );
  NAND2XL U1241 ( .A(n346), .B(n343), .Y(n129) );
  OR2X1 U1242 ( .A(n342), .B(n341), .Y(n982) );
  NAND2X1 U1243 ( .A(n342), .B(n341), .Y(n116) );
  INVX2 U1244 ( .A(n338), .Y(n339) );
  OR2X1 U1245 ( .A(n340), .B(n339), .Y(n983) );
  NAND2X1 U1246 ( .A(n340), .B(n339), .Y(n105) );
  NOR2X1 U1247 ( .A(n564), .B(n338), .Y(n91) );
  NAND2X1 U1248 ( .A(n564), .B(n338), .Y(n92) );
  ADDFHX1 U1249 ( .A(n616), .B(n661), .CI(n676), .CO(n446), .S(n447) );
  ADDFHX1 U1250 ( .A(n572), .B(n587), .CI(n602), .CO(n458), .S(n459) );
  ADDFHX1 U1251 ( .A(n556), .B(n617), .CI(n632), .CO(n460), .S(n461) );
  ADDFX1 U1252 ( .A(n573), .B(n678), .CI(n588), .CO(n474), .S(n475) );
  NOR2BXL U1253 ( .AN(b[0]), .B(n46), .Y(n573) );
  OAI2BB1X1 U1254 ( .A0N(n9), .A1N(n12), .B0(n554), .Y(n659) );
  ADDFHX1 U1255 ( .A(n646), .B(n586), .CI(n601), .CO(n444), .S(n445) );
  ADDHX1 U1256 ( .A(n677), .B(n647), .CO(n462), .S(n463) );
  OAI2BB1X1 U1257 ( .A0N(n34), .A1N(n36), .B0(n550), .Y(n591) );
  INVX2 U1258 ( .A(n726), .Y(n550) );
  ADDHX1 U1259 ( .A(n683), .B(n653), .CO(n522), .S(n523) );
  ADDFX1 U1260 ( .A(n624), .B(n684), .CI(n639), .CO(n528), .S(n529) );
  NOR2BXL U1261 ( .AN(b[0]), .B(n28), .Y(n624) );
  OAI22XL U1262 ( .A0(n12), .A1(n807), .B0(n806), .B1(n9), .Y(n672) );
  INVX2 U1263 ( .A(n988), .Y(n873) );
  OAI22XL U1264 ( .A0(n48), .A1(n701), .B0(n46), .B1(n700), .Y(n386) );
  OAI2BB1X1 U1265 ( .A0N(n954), .A1N(n24), .B0(n552), .Y(n625) );
  OAI22XL U1266 ( .A0(n12), .A1(n874), .B0(n9), .B1(n810), .Y(n562) );
  INVX2 U1267 ( .A(n987), .Y(n874) );
  OAI22XL U1268 ( .A0(n24), .A1(n959), .B0(n954), .B1(n776), .Y(n560) );
  NOR2BXL U1269 ( .AN(b[0]), .B(n40), .Y(n590) );
  ADDFX2 U1270 ( .A(n368), .B(n578), .CI(n608), .CO(n360), .S(n361) );
  OAI2BB1X1 U1271 ( .A0N(n28), .A1N(n30), .B0(n551), .Y(n608) );
  INVX2 U1272 ( .A(n743), .Y(n551) );
  INVX1 U1273 ( .A(n368), .Y(n369) );
  ADDFHX1 U1274 ( .A(n583), .B(n598), .CI(n628), .CO(n404), .S(n405) );
  XNOR2X1 U1275 ( .A(b[0]), .B(n986), .Y(n826) );
  NOR2BXL U1276 ( .AN(b[0]), .B(n34), .Y(n607) );
  INVX2 U1277 ( .A(n986), .Y(n875) );
  NAND2BX1 U1278 ( .AN(b[0]), .B(n986), .Y(n827) );
  ADDFHX1 U1279 ( .A(n569), .B(n582), .CI(n612), .CO(n394), .S(n395) );
  ADDFHX1 U1280 ( .A(n570), .B(n584), .CI(n644), .CO(n418), .S(n419) );
  INVX2 U1281 ( .A(n344), .Y(n345) );
  XNOR2X1 U1282 ( .A(b[0]), .B(n988), .Y(n792) );
  XNOR2X1 U1283 ( .A(b[0]), .B(n993), .Y(n707) );
  NAND2BX1 U1284 ( .AN(b[0]), .B(n993), .Y(n708) );
  XNOR2X1 U1285 ( .A(b[0]), .B(n987), .Y(n809) );
  XNOR2X1 U1286 ( .A(b[0]), .B(n991), .Y(n741) );
  NOR2BXL U1287 ( .AN(b[0]), .B(n9), .Y(n675) );
  XNOR2X1 U1288 ( .A(b[0]), .B(n990), .Y(n758) );
  NAND2BX1 U1289 ( .AN(b[0]), .B(n990), .Y(n759) );
  NAND2BX1 U1290 ( .AN(b[0]), .B(n987), .Y(n810) );
  INVX2 U1291 ( .A(n993), .Y(n868) );
  INVX2 U1292 ( .A(n991), .Y(n870) );
  INVX2 U1293 ( .A(n990), .Y(n871) );
  NOR2BXL U1294 ( .AN(b[0]), .B(n867), .Y(product[0]) );
  ADDFX2 U1295 ( .A(n344), .B(n565), .CI(n574), .CO(n340), .S(n341) );
  OAI2BB1X1 U1296 ( .A0N(n40), .A1N(n42), .B0(n549), .Y(n574) );
  INVX2 U1297 ( .A(n709), .Y(n549) );
  OAI2BB1X1 U1298 ( .A0N(n46), .A1N(n48), .B0(n548), .Y(n564) );
  INVX2 U1299 ( .A(n692), .Y(n548) );
  XOR2X1 U1300 ( .A(n987), .B(a[2]), .Y(n850) );
  XOR2X1 U1301 ( .A(n990), .B(a[8]), .Y(n847) );
  XNOR2X1 U1302 ( .A(n986), .B(b[14]), .Y(n812) );
  XOR2X2 U1303 ( .A(n986), .B(a[0]), .Y(n851) );
  XOR2X1 U1304 ( .A(n992), .B(a[12]), .Y(n845) );
  XNOR2X1 U1305 ( .A(n986), .B(b[13]), .Y(n813) );
  XNOR2X1 U1306 ( .A(n986), .B(b[15]), .Y(n811) );
  XNOR2X1 U1307 ( .A(n986), .B(b[10]), .Y(n816) );
  XNOR2X1 U1308 ( .A(n986), .B(b[8]), .Y(n818) );
  XNOR2X1 U1309 ( .A(n986), .B(b[7]), .Y(n819) );
  XNOR2X1 U1310 ( .A(n986), .B(b[4]), .Y(n822) );
  XNOR2X1 U1311 ( .A(n986), .B(b[12]), .Y(n814) );
  XNOR2X1 U1312 ( .A(n986), .B(b[9]), .Y(n817) );
  XNOR2X1 U1313 ( .A(n986), .B(b[2]), .Y(n824) );
  XNOR2X1 U1314 ( .A(n986), .B(b[1]), .Y(n825) );
  XNOR2X1 U1315 ( .A(n986), .B(b[3]), .Y(n823) );
  XNOR2X1 U1316 ( .A(n988), .B(b[15]), .Y(n777) );
  XNOR2X1 U1317 ( .A(n990), .B(b[6]), .Y(n752) );
  XNOR2X1 U1318 ( .A(n987), .B(b[15]), .Y(n794) );
  XNOR2X1 U1319 ( .A(n988), .B(b[7]), .Y(n785) );
  XNOR2X1 U1320 ( .A(n988), .B(b[12]), .Y(n780) );
  XNOR2X1 U1321 ( .A(n988), .B(b[4]), .Y(n788) );
  XNOR2X1 U1322 ( .A(n987), .B(b[12]), .Y(n797) );
  XNOR2X1 U1323 ( .A(n988), .B(b[5]), .Y(n787) );
  XNOR2X1 U1324 ( .A(n992), .B(b[3]), .Y(n721) );
  XNOR2X1 U1325 ( .A(n990), .B(b[5]), .Y(n753) );
  XNOR2X1 U1326 ( .A(n990), .B(b[7]), .Y(n751) );
  XNOR2X1 U1327 ( .A(n987), .B(b[13]), .Y(n796) );
  XNOR2X1 U1328 ( .A(n988), .B(b[11]), .Y(n781) );
  XNOR2X1 U1329 ( .A(n988), .B(b[3]), .Y(n789) );
  XNOR2X1 U1330 ( .A(n988), .B(b[14]), .Y(n778) );
  XNOR2X1 U1331 ( .A(n992), .B(b[4]), .Y(n720) );
  XNOR2X1 U1332 ( .A(n992), .B(b[2]), .Y(n722) );
  XNOR2X1 U1333 ( .A(n990), .B(b[8]), .Y(n750) );
  XNOR2X1 U1334 ( .A(n988), .B(b[13]), .Y(n779) );
  XNOR2X1 U1335 ( .A(n989), .B(b[10]), .Y(n765) );
  XNOR2X1 U1336 ( .A(n987), .B(b[10]), .Y(n799) );
  XNOR2X1 U1337 ( .A(n991), .B(b[4]), .Y(n737) );
  XNOR2X1 U1338 ( .A(n990), .B(b[9]), .Y(n749) );
  XNOR2X1 U1339 ( .A(n991), .B(b[8]), .Y(n733) );
  XNOR2X1 U1340 ( .A(n988), .B(b[10]), .Y(n782) );
  XNOR2X1 U1341 ( .A(n989), .B(b[8]), .Y(n767) );
  XNOR2X1 U1342 ( .A(n989), .B(b[4]), .Y(n771) );
  XNOR2X1 U1343 ( .A(n988), .B(b[9]), .Y(n783) );
  XNOR2X1 U1344 ( .A(n987), .B(b[9]), .Y(n800) );
  XNOR2X1 U1345 ( .A(n992), .B(b[1]), .Y(n723) );
  XNOR2X1 U1346 ( .A(n989), .B(b[9]), .Y(n766) );
  XNOR2X1 U1347 ( .A(n991), .B(b[1]), .Y(n740) );
  XNOR2X1 U1348 ( .A(n991), .B(b[3]), .Y(n738) );
  XNOR2X1 U1349 ( .A(n991), .B(b[7]), .Y(n734) );
  XNOR2X1 U1350 ( .A(n992), .B(b[5]), .Y(n719) );
  XNOR2X1 U1351 ( .A(n989), .B(b[7]), .Y(n768) );
  XNOR2X1 U1352 ( .A(n989), .B(b[3]), .Y(n772) );
  XNOR2X1 U1353 ( .A(n990), .B(b[3]), .Y(n755) );
  XNOR2X1 U1354 ( .A(n988), .B(b[1]), .Y(n791) );
  XNOR2X1 U1355 ( .A(n989), .B(b[6]), .Y(n769) );
  XNOR2X1 U1356 ( .A(n988), .B(b[8]), .Y(n784) );
  XNOR2X1 U1357 ( .A(n989), .B(b[5]), .Y(n770) );
  XNOR2X1 U1358 ( .A(n988), .B(b[2]), .Y(n790) );
  XNOR2X1 U1359 ( .A(n990), .B(b[1]), .Y(n757) );
  XNOR2X1 U1360 ( .A(n991), .B(b[2]), .Y(n739) );
  XNOR2X1 U1361 ( .A(n991), .B(b[9]), .Y(n732) );
  XNOR2X1 U1362 ( .A(n987), .B(b[2]), .Y(n807) );
  XNOR2X1 U1363 ( .A(n990), .B(b[2]), .Y(n756) );
  XNOR2X1 U1364 ( .A(n990), .B(b[10]), .Y(n748) );
  XNOR2X1 U1365 ( .A(n992), .B(b[7]), .Y(n717) );
  XNOR2X1 U1366 ( .A(n989), .B(b[1]), .Y(n774) );
  XNOR2X1 U1367 ( .A(n992), .B(b[8]), .Y(n716) );
  XNOR2X1 U1368 ( .A(n992), .B(b[6]), .Y(n718) );
  XNOR2X1 U1369 ( .A(n992), .B(b[10]), .Y(n714) );
  XNOR2X1 U1370 ( .A(n989), .B(b[15]), .Y(n760) );
  XNOR2X1 U1371 ( .A(n987), .B(b[6]), .Y(n803) );
  XNOR2X1 U1372 ( .A(n990), .B(b[4]), .Y(n754) );
  XNOR2X1 U1373 ( .A(n987), .B(b[1]), .Y(n808) );
  XNOR2X1 U1374 ( .A(n987), .B(b[3]), .Y(n806) );
  XNOR2X1 U1375 ( .A(n991), .B(b[10]), .Y(n731) );
  XNOR2X1 U1376 ( .A(n989), .B(b[2]), .Y(n773) );
  XNOR2X1 U1377 ( .A(n992), .B(b[9]), .Y(n715) );
  XNOR2X1 U1378 ( .A(n987), .B(b[5]), .Y(n804) );
  XNOR2X1 U1379 ( .A(n991), .B(b[11]), .Y(n730) );
  XNOR2X1 U1380 ( .A(n987), .B(b[8]), .Y(n801) );
  XNOR2X1 U1381 ( .A(n991), .B(b[12]), .Y(n729) );
  XNOR2X1 U1382 ( .A(n992), .B(b[11]), .Y(n713) );
  XNOR2X1 U1383 ( .A(n991), .B(b[13]), .Y(n728) );
  XNOR2X1 U1384 ( .A(n989), .B(b[14]), .Y(n761) );
  XNOR2X1 U1385 ( .A(n991), .B(b[5]), .Y(n736) );
  XNOR2X1 U1386 ( .A(n987), .B(b[4]), .Y(n805) );
  XNOR2X1 U1387 ( .A(n992), .B(b[13]), .Y(n711) );
  XNOR2X1 U1388 ( .A(n991), .B(b[6]), .Y(n735) );
  XNOR2X1 U1389 ( .A(n992), .B(b[14]), .Y(n710) );
  XNOR2X1 U1390 ( .A(n992), .B(b[12]), .Y(n712) );
  XNOR2X1 U1391 ( .A(n987), .B(b[7]), .Y(n802) );
  XNOR2X1 U1392 ( .A(n989), .B(b[12]), .Y(n763) );
  XNOR2X1 U1393 ( .A(n989), .B(b[11]), .Y(n764) );
  XNOR2X1 U1394 ( .A(n990), .B(b[12]), .Y(n746) );
  XNOR2X1 U1395 ( .A(n989), .B(b[13]), .Y(n762) );
  XNOR2X1 U1396 ( .A(n991), .B(b[14]), .Y(n727) );
  XNOR2X1 U1397 ( .A(n990), .B(b[13]), .Y(n745) );
  XNOR2X1 U1398 ( .A(n990), .B(b[15]), .Y(n743) );
  BUFX2 U1399 ( .A(n664), .Y(n984) );
  OAI22XL U1400 ( .A0(n12), .A1(n799), .B0(n798), .B1(n9), .Y(n664) );
  ADDHXL U1401 ( .A(n685), .B(n655), .CO(n534), .S(n535) );
  OAI22XL U1402 ( .A0(n12), .A1(n798), .B0(n797), .B1(n9), .Y(n663) );
  OAI2BB1X1 U1403 ( .A0N(n867), .A1N(n6), .B0(n555), .Y(n676) );
  OAI22XL U1404 ( .A0(n6), .A1(n814), .B0(n813), .B1(n867), .Y(n679) );
  OAI22XL U1405 ( .A0(n6), .A1(n813), .B0(n812), .B1(n867), .Y(n678) );
  OAI22XL U1406 ( .A0(n6), .A1(n875), .B0(n827), .B1(n867), .Y(n563) );
  OAI22XL U1407 ( .A0(n6), .A1(n821), .B0(n820), .B1(n867), .Y(n686) );
  OAI22XL U1408 ( .A0(n6), .A1(n825), .B0(n824), .B1(n867), .Y(n690) );
  OAI22XL U1409 ( .A0(n826), .A1(n6), .B0(n825), .B1(n867), .Y(n691) );
  OAI22XL U1410 ( .A0(n18), .A1(n779), .B0(n778), .B1(n951), .Y(n644) );
  OAI2BB1X1 U1411 ( .A0N(n951), .A1N(n18), .B0(n553), .Y(n642) );
  OAI22XL U1412 ( .A0(n18), .A1(n785), .B0(n784), .B1(n951), .Y(n650) );
  OAI22XL U1413 ( .A0(n18), .A1(n783), .B0(n782), .B1(n951), .Y(n648) );
  OAI22XL U1414 ( .A0(n18), .A1(n780), .B0(n779), .B1(n951), .Y(n645) );
  OAI22XL U1415 ( .A0(n18), .A1(n791), .B0(n790), .B1(n951), .Y(n656) );
  OAI22XL U1416 ( .A0(n18), .A1(n789), .B0(n788), .B1(n951), .Y(n654) );
  NOR2BXL U1417 ( .AN(b[0]), .B(n951), .Y(n658) );
  OAI22XL U1418 ( .A0(n18), .A1(n873), .B0(n951), .B1(n793), .Y(n561) );
  OAI22XL U1419 ( .A0(n18), .A1(n790), .B0(n789), .B1(n951), .Y(n655) );
  OAI22XL U1420 ( .A0(n18), .A1(n781), .B0(n780), .B1(n951), .Y(n646) );
  ADDHXL U1421 ( .A(n679), .B(n649), .CO(n486), .S(n487) );
  OAI22XL U1422 ( .A0(n18), .A1(n784), .B0(n783), .B1(n951), .Y(n649) );
  NOR2X4 U1423 ( .A(n437), .B(n450), .Y(n227) );
  OAI21XL U1424 ( .A0(n211), .A1(n219), .B0(n212), .Y(n210) );
  XOR2X2 U1425 ( .A(n130), .B(n57), .Y(product[27]) );
  OAI22X2 U1426 ( .A0(n48), .A1(n705), .B0(n46), .B1(n704), .Y(n434) );
  OAI21XL U1427 ( .A0(n224), .A1(n216), .B0(n219), .Y(n215) );
  OR2X1 U1428 ( .A(n631), .B(n571), .Y(n448) );
  XOR2X2 U1429 ( .A(n106), .B(n55), .Y(product[29]) );
  AOI21X4 U1430 ( .A0(n255), .A1(n236), .B0(n237), .Y(n235) );
endmodule


module PE_DW01_add_26 ( A, B, CI, SUM, CO );
  input [36:0] A;
  input [36:0] B;
  output [36:0] SUM;
  input CI;
  output CO;
  wire   n3, n4, n6, n8, n9, n10, n11, n13, n15, n16, n17, n18, n19, n20, n21,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n56, n57, n58, n59, n60, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n87, n89, n90,
         n91, n92, n94, n97, n98, n99, n100, n101, n103, n105, n108, n109,
         n110, n111, n113, n115, n116, n117, n118, n119, n120, n121, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n140, n142, n143, n145, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n162, n164, n165, n167, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n197, n199,
         n200, n201, n202, n203, n205, n207, n208, n209, n210, n211, n213,
         n214, n215, n216, n218, n219, n220, n221, n230, n231, n233, n236,
         n237, n240, n241, n242, n243, n244, n245, n250, n252, n253, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395;

  OAI21X4 U11 ( .A0(n42), .A1(n40), .B0(n41), .Y(n39) );
  NAND2X4 U15 ( .A(B[31]), .B(A[31]), .Y(n41) );
  AOI21X1 U73 ( .A0(n94), .A1(n372), .B0(n87), .Y(n83) );
  XNOR2X4 U82 ( .A(n101), .B(n10), .Y(SUM[24]) );
  AOI21X1 U118 ( .A0(n126), .A1(n117), .B0(n118), .Y(n116) );
  NOR2X2 U131 ( .A(A[20]), .B(B[20]), .Y(n124) );
  OAI21X4 U150 ( .A0(n149), .A1(n137), .B0(n138), .Y(n136) );
  XNOR2X4 U291 ( .A(n39), .B(n385), .Y(SUM[32]) );
  XNOR2X2 U292 ( .A(n132), .B(n15), .Y(SUM[19]) );
  NAND2X2 U293 ( .A(A[14]), .B(B[14]), .Y(n156) );
  NOR2X1 U294 ( .A(A[15]), .B(B[15]), .Y(n152) );
  NOR2X2 U295 ( .A(A[19]), .B(B[19]), .Y(n130) );
  OAI21X1 U296 ( .A0(n179), .A1(n177), .B0(n178), .Y(n176) );
  OAI21X1 U297 ( .A0(n92), .A1(n75), .B0(n76), .Y(n74) );
  AOI21X4 U298 ( .A0(n388), .A1(n145), .B0(n140), .Y(n138) );
  XOR2X2 U299 ( .A(n50), .B(n4), .Y(SUM[30]) );
  NAND2XL U300 ( .A(A[22]), .B(B[22]), .Y(n115) );
  INVX3 U301 ( .A(n72), .Y(n71) );
  NAND2X2 U302 ( .A(n380), .B(n103), .Y(n101) );
  AOI21X2 U303 ( .A0(n77), .A1(n87), .B0(n78), .Y(n76) );
  NOR2X2 U304 ( .A(B[11]), .B(A[11]), .Y(n174) );
  XOR2X2 U305 ( .A(n57), .B(n384), .Y(SUM[29]) );
  NAND2X2 U306 ( .A(n361), .B(n362), .Y(n363) );
  NAND2X2 U307 ( .A(n363), .B(n65), .Y(n59) );
  INVX1 U308 ( .A(n64), .Y(n361) );
  INVX2 U309 ( .A(n70), .Y(n362) );
  NOR2X2 U310 ( .A(A[28]), .B(B[28]), .Y(n64) );
  OAI2BB1X2 U311 ( .A0N(n59), .A1N(n374), .B0(n56), .Y(n52) );
  AOI21X1 U312 ( .A0(n46), .A1(n59), .B0(n47), .Y(n45) );
  NAND2XL U313 ( .A(n71), .B(n67), .Y(n364) );
  INVX2 U314 ( .A(n68), .Y(n365) );
  AND2X4 U315 ( .A(n364), .B(n365), .Y(n66) );
  XOR2X4 U316 ( .A(n66), .B(n6), .Y(SUM[28]) );
  NAND2X2 U317 ( .A(n366), .B(n367), .Y(n368) );
  NAND2X2 U318 ( .A(n368), .B(n45), .Y(n43) );
  CLKINVX2 U319 ( .A(n72), .Y(n366) );
  CLKINVX2 U320 ( .A(n44), .Y(n367) );
  AOI21X1 U321 ( .A0(n43), .A1(n35), .B0(n36), .Y(SUM[34]) );
  INVX4 U322 ( .A(n43), .Y(n42) );
  AOI21X1 U323 ( .A0(n71), .A1(n58), .B0(n59), .Y(n57) );
  NAND2X1 U324 ( .A(n117), .B(n371), .Y(n110) );
  NAND2XL U325 ( .A(n58), .B(n46), .Y(n44) );
  XNOR2X2 U326 ( .A(n81), .B(n8), .Y(SUM[26]) );
  XOR2X1 U327 ( .A(n387), .B(n216), .Y(SUM[1]) );
  NAND2XL U328 ( .A(n221), .B(n49), .Y(n4) );
  OAI21X2 U329 ( .A0(n127), .A1(n110), .B0(n111), .Y(n109) );
  NAND2XL U330 ( .A(n392), .B(n391), .Y(n159) );
  NOR2X1 U331 ( .A(A[6]), .B(B[6]), .Y(n193) );
  OAI21X1 U332 ( .A0(n193), .A1(n195), .B0(n194), .Y(n192) );
  NAND2X1 U333 ( .A(A[20]), .B(B[20]), .Y(n125) );
  XNOR2X1 U334 ( .A(n31), .B(n208), .Y(SUM[3]) );
  XOR2X1 U335 ( .A(n30), .B(n203), .Y(SUM[4]) );
  NAND2X1 U336 ( .A(A[7]), .B(B[7]), .Y(n190) );
  NOR2X2 U337 ( .A(A[21]), .B(B[21]), .Y(n119) );
  NAND2X1 U338 ( .A(A[21]), .B(B[21]), .Y(n120) );
  OR2X2 U339 ( .A(n378), .B(n94), .Y(n90) );
  AOI21X2 U340 ( .A0(n109), .A1(n73), .B0(n74), .Y(n72) );
  NOR2X1 U341 ( .A(n91), .B(n75), .Y(n73) );
  INVX1 U342 ( .A(A[33]), .Y(n253) );
  INVX1 U343 ( .A(B[33]), .Y(n252) );
  OAI21X1 U344 ( .A0(n183), .A1(n181), .B0(n182), .Y(n180) );
  NOR2X1 U345 ( .A(A[1]), .B(B[1]), .Y(n214) );
  OAI21X1 U346 ( .A0(n211), .A1(n209), .B0(n210), .Y(n208) );
  NOR2X1 U347 ( .A(A[4]), .B(B[4]), .Y(n201) );
  AOI21X2 U348 ( .A0(n150), .A1(n158), .B0(n151), .Y(n149) );
  OAI21X1 U349 ( .A0(n152), .A1(n156), .B0(n153), .Y(n151) );
  NOR2X1 U350 ( .A(n155), .B(n152), .Y(n150) );
  NOR2X1 U351 ( .A(n60), .B(n53), .Y(n51) );
  NAND2X1 U352 ( .A(A[24]), .B(B[24]), .Y(n100) );
  NOR2X2 U353 ( .A(A[24]), .B(B[24]), .Y(n99) );
  NOR2X1 U354 ( .A(A[2]), .B(B[2]), .Y(n209) );
  NAND2X1 U355 ( .A(n245), .B(n194), .Y(n28) );
  XOR2X1 U356 ( .A(n165), .B(n21), .Y(SUM[13]) );
  OR2X1 U357 ( .A(n376), .B(n377), .Y(n132) );
  XNOR2X1 U358 ( .A(n154), .B(n19), .Y(SUM[15]) );
  OR2X1 U359 ( .A(A[16]), .B(B[16]), .Y(n389) );
  NOR2X1 U360 ( .A(n124), .B(n119), .Y(n117) );
  NAND2X2 U361 ( .A(A[23]), .B(B[23]), .Y(n103) );
  NOR2X1 U362 ( .A(A[27]), .B(B[27]), .Y(n69) );
  NAND2X1 U363 ( .A(A[27]), .B(B[27]), .Y(n70) );
  XNOR2X1 U364 ( .A(n26), .B(n188), .Y(SUM[8]) );
  NAND2X1 U365 ( .A(n243), .B(n187), .Y(n26) );
  OAI21X1 U366 ( .A0(n375), .A1(n191), .B0(n190), .Y(n188) );
  OAI21X1 U367 ( .A0(n108), .A1(n82), .B0(n83), .Y(n81) );
  XOR2X1 U368 ( .A(n121), .B(n13), .Y(SUM[21]) );
  NAND2X1 U369 ( .A(n230), .B(n120), .Y(n13) );
  NOR2X1 U370 ( .A(n69), .B(n64), .Y(n58) );
  NOR2X1 U371 ( .A(n48), .B(n53), .Y(n46) );
  NOR2X1 U372 ( .A(B[30]), .B(A[30]), .Y(n48) );
  NAND2X1 U373 ( .A(B[30]), .B(A[30]), .Y(n49) );
  NOR2X1 U374 ( .A(n40), .B(n37), .Y(n35) );
  OAI21X2 U375 ( .A0(n171), .A1(n159), .B0(n160), .Y(n158) );
  OR2X4 U376 ( .A(B[23]), .B(A[23]), .Y(n369) );
  AND2X1 U377 ( .A(n373), .B(n218), .Y(SUM[0]) );
  AOI21X1 U378 ( .A0(n172), .A1(n180), .B0(n173), .Y(n171) );
  OR2X4 U379 ( .A(A[22]), .B(B[22]), .Y(n371) );
  OR2X4 U380 ( .A(A[25]), .B(B[25]), .Y(n372) );
  OR2X1 U381 ( .A(A[0]), .B(B[0]), .Y(n373) );
  AOI21X1 U382 ( .A0(n184), .A1(n192), .B0(n185), .Y(n183) );
  NAND2X2 U383 ( .A(n388), .B(n389), .Y(n137) );
  INVX2 U384 ( .A(n127), .Y(n126) );
  AOI21X2 U385 ( .A0(n392), .A1(n167), .B0(n162), .Y(n160) );
  XNOR2X1 U386 ( .A(n116), .B(n390), .Y(SUM[22]) );
  NAND2X4 U387 ( .A(n372), .B(n77), .Y(n75) );
  INVX3 U388 ( .A(n109), .Y(n108) );
  OR2X1 U389 ( .A(A[29]), .B(B[29]), .Y(n374) );
  INVX1 U390 ( .A(n244), .Y(n375) );
  CLKINVXL U391 ( .A(n189), .Y(n244) );
  NOR2X1 U392 ( .A(n135), .B(n133), .Y(n376) );
  CLKINVXL U393 ( .A(n134), .Y(n377) );
  NOR2X1 U394 ( .A(B[18]), .B(A[18]), .Y(n133) );
  NAND2X1 U395 ( .A(B[18]), .B(A[18]), .Y(n134) );
  NAND2X4 U396 ( .A(n369), .B(n97), .Y(n91) );
  NAND2XL U397 ( .A(A[28]), .B(B[28]), .Y(n65) );
  INVX1 U398 ( .A(n214), .Y(n250) );
  NOR2X1 U399 ( .A(n108), .B(n91), .Y(n378) );
  OAI21X2 U400 ( .A0(n130), .A1(n134), .B0(n131), .Y(n129) );
  CLKINVXL U401 ( .A(n108), .Y(n379) );
  NAND2X1 U402 ( .A(n253), .B(n252), .Y(n38) );
  XOR2X1 U403 ( .A(n170), .B(n386), .Y(SUM[12]) );
  NOR2X2 U404 ( .A(n253), .B(n252), .Y(n37) );
  NAND2X1 U405 ( .A(n379), .B(n369), .Y(n380) );
  NOR2X2 U406 ( .A(n130), .B(n133), .Y(n128) );
  INVX1 U407 ( .A(n180), .Y(n179) );
  NAND2BX1 U408 ( .AN(n130), .B(n131), .Y(n15) );
  NAND2XL U409 ( .A(A[16]), .B(B[16]), .Y(n147) );
  INVX2 U410 ( .A(n192), .Y(n191) );
  NAND2XL U411 ( .A(n374), .B(n56), .Y(n384) );
  NOR2X1 U412 ( .A(A[7]), .B(B[7]), .Y(n189) );
  CLKINVXL U413 ( .A(n133), .Y(n233) );
  AOI21XL U414 ( .A0(n148), .A1(n389), .B0(n145), .Y(n143) );
  INVX4 U415 ( .A(n103), .Y(n105) );
  INVX3 U416 ( .A(n100), .Y(n98) );
  AND2X1 U417 ( .A(n240), .B(n175), .Y(n382) );
  NAND2X1 U418 ( .A(n242), .B(n182), .Y(n25) );
  OAI21XL U419 ( .A0(n48), .A1(n56), .B0(n49), .Y(n47) );
  INVX1 U420 ( .A(n164), .Y(n162) );
  NAND2XL U421 ( .A(n392), .B(n164), .Y(n21) );
  XNOR2X1 U422 ( .A(n71), .B(n383), .Y(SUM[27]) );
  NAND2XL U423 ( .A(n67), .B(n70), .Y(n383) );
  INVX1 U424 ( .A(n199), .Y(n197) );
  CLKINVXL U425 ( .A(n69), .Y(n67) );
  OR2X4 U426 ( .A(A[13]), .B(B[13]), .Y(n392) );
  INVX3 U427 ( .A(n79), .Y(n77) );
  NAND2XL U428 ( .A(A[2]), .B(B[2]), .Y(n210) );
  NAND2X1 U429 ( .A(A[1]), .B(B[1]), .Y(n215) );
  CLKINVXL U430 ( .A(n136), .Y(n135) );
  XOR2X1 U431 ( .A(n135), .B(n16), .Y(SUM[18]) );
  XOR2X1 U432 ( .A(n143), .B(n17), .Y(SUM[17]) );
  XOR2X1 U433 ( .A(n126), .B(n381), .Y(SUM[20]) );
  AND2X1 U434 ( .A(n231), .B(n125), .Y(n381) );
  XNOR2X1 U435 ( .A(n148), .B(n18), .Y(SUM[16]) );
  CLKINVXL U436 ( .A(n171), .Y(n170) );
  OR2X4 U437 ( .A(A[17]), .B(B[17]), .Y(n388) );
  NAND2XL U438 ( .A(n97), .B(n100), .Y(n10) );
  NAND2XL U439 ( .A(A[17]), .B(B[17]), .Y(n142) );
  XOR2X1 U440 ( .A(n157), .B(n20), .Y(SUM[14]) );
  CLKINVXL U441 ( .A(n155), .Y(n237) );
  NAND2XL U442 ( .A(n236), .B(n153), .Y(n19) );
  OAI21XL U443 ( .A0(n157), .A1(n155), .B0(n156), .Y(n154) );
  XOR2X1 U444 ( .A(n176), .B(n382), .Y(SUM[11]) );
  XOR2XL U445 ( .A(n24), .B(n179), .Y(SUM[10]) );
  NAND2XL U446 ( .A(n241), .B(n178), .Y(n24) );
  CLKINVXL U447 ( .A(n177), .Y(n241) );
  XOR2XL U448 ( .A(n25), .B(n183), .Y(SUM[9]) );
  CLKINVXL U449 ( .A(n181), .Y(n242) );
  AOI21X1 U450 ( .A0(n71), .A1(n51), .B0(n52), .Y(n50) );
  NAND2X4 U451 ( .A(n220), .B(n41), .Y(n3) );
  XOR2X4 U452 ( .A(n42), .B(n3), .Y(SUM[31]) );
  NAND2BX1 U453 ( .AN(n64), .B(n65), .Y(n6) );
  INVX1 U454 ( .A(n169), .Y(n167) );
  NAND2X4 U455 ( .A(n219), .B(n38), .Y(n385) );
  OAI21X1 U456 ( .A0(n186), .A1(n190), .B0(n187), .Y(n185) );
  AOI21X1 U457 ( .A0(n394), .A1(n200), .B0(n197), .Y(n195) );
  AND2X1 U458 ( .A(n391), .B(n169), .Y(n386) );
  AOI21XL U459 ( .A0(n170), .A1(n391), .B0(n167), .Y(n165) );
  XOR2X1 U460 ( .A(n27), .B(n191), .Y(SUM[7]) );
  XNOR2XL U461 ( .A(n29), .B(n200), .Y(SUM[5]) );
  NAND2XL U462 ( .A(n394), .B(n199), .Y(n29) );
  CLKINVXL U463 ( .A(n193), .Y(n245) );
  XOR2XL U464 ( .A(n28), .B(n195), .Y(SUM[6]) );
  NAND2BX1 U465 ( .AN(n201), .B(n202), .Y(n30) );
  NAND2XL U466 ( .A(A[13]), .B(B[13]), .Y(n164) );
  OR2X2 U467 ( .A(A[3]), .B(B[3]), .Y(n393) );
  NAND2XL U468 ( .A(A[3]), .B(B[3]), .Y(n207) );
  NAND2X1 U469 ( .A(A[6]), .B(B[6]), .Y(n194) );
  NAND2XL U470 ( .A(A[4]), .B(B[4]), .Y(n202) );
  OR2X2 U471 ( .A(A[5]), .B(B[5]), .Y(n394) );
  NAND2BX1 U472 ( .AN(n209), .B(n210), .Y(n32) );
  AND2X1 U473 ( .A(n250), .B(n215), .Y(n387) );
  INVX2 U474 ( .A(n142), .Y(n140) );
  NAND2X1 U475 ( .A(n388), .B(n142), .Y(n17) );
  INVX2 U476 ( .A(n147), .Y(n145) );
  NAND2X1 U477 ( .A(n233), .B(n134), .Y(n16) );
  INVX2 U478 ( .A(n124), .Y(n231) );
  CLKINVXL U479 ( .A(n125), .Y(n123) );
  INVX2 U480 ( .A(n395), .Y(SUM[35]) );
  INVX2 U481 ( .A(n395), .Y(SUM[36]) );
  INVX2 U482 ( .A(n395), .Y(SUM[33]) );
  INVX2 U483 ( .A(n115), .Y(n113) );
  NAND2XL U484 ( .A(n372), .B(n89), .Y(n9) );
  INVXL U485 ( .A(n174), .Y(n240) );
  OAI21X1 U486 ( .A0(n174), .A1(n178), .B0(n175), .Y(n173) );
  CLKINVXL U487 ( .A(n119), .Y(n230) );
  CLKINVXL U488 ( .A(n158), .Y(n157) );
  CLKINVXL U489 ( .A(n152), .Y(n236) );
  AND2X1 U490 ( .A(n371), .B(n115), .Y(n390) );
  NAND2BX1 U491 ( .AN(n91), .B(n372), .Y(n82) );
  NAND2X1 U492 ( .A(A[19]), .B(B[19]), .Y(n131) );
  NAND2XL U493 ( .A(n237), .B(n156), .Y(n20) );
  CLKINVXL U494 ( .A(SUM[34]), .Y(n395) );
  CLKINVXL U495 ( .A(n48), .Y(n221) );
  OAI21XL U496 ( .A0(n41), .A1(n37), .B0(n38), .Y(n36) );
  NOR2X1 U497 ( .A(B[9]), .B(A[9]), .Y(n181) );
  NOR2X1 U498 ( .A(n186), .B(n189), .Y(n184) );
  NOR2X1 U499 ( .A(B[8]), .B(A[8]), .Y(n186) );
  NOR2X1 U500 ( .A(B[10]), .B(A[10]), .Y(n177) );
  NOR2X1 U501 ( .A(A[14]), .B(B[14]), .Y(n155) );
  OAI21XL U502 ( .A0(n203), .A1(n201), .B0(n202), .Y(n200) );
  CLKINVXL U503 ( .A(n186), .Y(n243) );
  NAND2X1 U504 ( .A(B[8]), .B(A[8]), .Y(n187) );
  NAND2X1 U505 ( .A(B[10]), .B(A[10]), .Y(n178) );
  NAND2X1 U506 ( .A(B[11]), .B(A[11]), .Y(n175) );
  NAND2XL U507 ( .A(n244), .B(n190), .Y(n27) );
  AOI21X1 U508 ( .A0(n208), .A1(n393), .B0(n205), .Y(n203) );
  INVX2 U509 ( .A(n207), .Y(n205) );
  NAND2X1 U510 ( .A(B[9]), .B(A[9]), .Y(n182) );
  NAND2X1 U511 ( .A(A[15]), .B(B[15]), .Y(n153) );
  NAND2X1 U512 ( .A(n393), .B(n207), .Y(n31) );
  CLKINVXL U513 ( .A(n70), .Y(n68) );
  NOR2X1 U514 ( .A(A[29]), .B(B[29]), .Y(n53) );
  NAND2X1 U515 ( .A(A[29]), .B(B[29]), .Y(n56) );
  OR2X1 U516 ( .A(A[12]), .B(B[12]), .Y(n391) );
  NAND2X1 U517 ( .A(A[12]), .B(B[12]), .Y(n169) );
  NAND2X1 U518 ( .A(A[5]), .B(B[5]), .Y(n199) );
  AOI21X1 U519 ( .A0(n250), .A1(n216), .B0(n213), .Y(n211) );
  INVX2 U520 ( .A(n215), .Y(n213) );
  INVX2 U521 ( .A(n218), .Y(n216) );
  NAND2X1 U522 ( .A(A[0]), .B(B[0]), .Y(n218) );
  CLKINVXL U523 ( .A(n92), .Y(n94) );
  INVX1 U524 ( .A(n80), .Y(n78) );
  NAND2XL U525 ( .A(n77), .B(n80), .Y(n8) );
  NAND2X1 U526 ( .A(B[26]), .B(A[26]), .Y(n80) );
  CLKINVX2 U527 ( .A(n149), .Y(n148) );
  CLKINVXL U528 ( .A(n58), .Y(n60) );
  AOI21X4 U529 ( .A0(n128), .A1(n136), .B0(n129), .Y(n127) );
  NAND2XL U530 ( .A(n389), .B(n147), .Y(n18) );
  XOR2X2 U531 ( .A(n108), .B(n11), .Y(SUM[23]) );
  AOI21X2 U532 ( .A0(n118), .A1(n371), .B0(n113), .Y(n111) );
  INVX4 U533 ( .A(n99), .Y(n97) );
  NAND2XL U534 ( .A(n369), .B(n103), .Y(n11) );
  OAI21X2 U535 ( .A0(n119), .A1(n125), .B0(n120), .Y(n118) );
  NOR2X4 U536 ( .A(A[26]), .B(B[26]), .Y(n79) );
  INVX2 U537 ( .A(n40), .Y(n220) );
  NOR2X4 U538 ( .A(B[31]), .B(A[31]), .Y(n40) );
  NAND2X2 U539 ( .A(A[25]), .B(B[25]), .Y(n89) );
  INVX2 U540 ( .A(n89), .Y(n87) );
  AOI21X4 U541 ( .A0(n97), .A1(n105), .B0(n98), .Y(n92) );
  XNOR2X4 U542 ( .A(n90), .B(n9), .Y(SUM[25]) );
  AOI21X2 U543 ( .A0(n126), .A1(n231), .B0(n123), .Y(n121) );
  NOR2X1 U544 ( .A(n177), .B(n174), .Y(n172) );
  XOR2X1 U545 ( .A(n32), .B(n211), .Y(SUM[2]) );
  CLKINVX8 U546 ( .A(n37), .Y(n219) );
endmodule


module PE_DW01_add_24 ( A, B, CI, SUM, CO );
  input [35:0] A;
  input [35:0] B;
  output [35:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n7, n9, n10, n11, n13, n14, n15, n16, n17, n20, n21, n22,
         n24, n25, n26, n28, n29, n30, n31, n32, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n50, n51, n52, n53, n54, n55, n57,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n115, n116, n117, n118,
         n120, n123, n124, n125, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n137, n139, n140, n141, n142, n146, n147, n148, n149,
         n150, n151, n152, n153, n157, n159, n160, n161, n162, n164, n167,
         n168, n169, n170, n172, n174, n175, n177, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n196,
         n197, n199, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n217, n219, n220, n221, n222,
         n223, n225, n227, n228, n229, n230, n231, n233, n235, n236, n237,
         n238, n240, n242, n243, n245, n247, n248, n250, n251, n252, n254,
         n256, n259, n260, n263, n265, n267, n269, n271, n273, n274, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411;

  AOI21X1 U7 ( .A0(n55), .A1(n38), .B0(n39), .Y(n37) );
  AOI21X1 U29 ( .A0(n73), .A1(n54), .B0(n55), .Y(n53) );
  AOI21X1 U43 ( .A0(n73), .A1(n65), .B0(n66), .Y(n64) );
  XNOR2X4 U64 ( .A(n87), .B(n7), .Y(SUM[26]) );
  OAI21X4 U75 ( .A0(n101), .A1(n88), .B0(n89), .Y(n87) );
  OAI21X4 U89 ( .A0(n101), .A1(n99), .B0(n100), .Y(n98) );
  AOI21X1 U116 ( .A0(n130), .A1(n117), .B0(n118), .Y(n116) );
  AOI21X1 U141 ( .A0(n405), .A1(n146), .B0(n137), .Y(n135) );
  AOI21X1 U151 ( .A0(n153), .A1(n254), .B0(n146), .Y(n142) );
  AOI21X1 U188 ( .A0(n406), .A1(n177), .B0(n172), .Y(n170) );
  XOR2X4 U311 ( .A(n125), .B(n394), .Y(SUM[21]) );
  AOI21X2 U312 ( .A0(n180), .A1(n407), .B0(n177), .Y(n175) );
  INVX2 U313 ( .A(n181), .Y(n180) );
  XOR2X2 U314 ( .A(n175), .B(n393), .Y(SUM[15]) );
  INVX2 U315 ( .A(n203), .Y(n202) );
  AOI21X4 U316 ( .A0(n130), .A1(n252), .B0(n127), .Y(n125) );
  INVX4 U317 ( .A(n131), .Y(n130) );
  XNOR2X2 U318 ( .A(n62), .B(n4), .Y(SUM[29]) );
  AND2X4 U319 ( .A(n390), .B(n164), .Y(n379) );
  NOR2X4 U320 ( .A(n379), .B(n157), .Y(n151) );
  OR2X2 U321 ( .A(A[17]), .B(B[17]), .Y(n390) );
  INVX20 U322 ( .A(n159), .Y(n157) );
  INVX1 U323 ( .A(n151), .Y(n153) );
  NAND2X2 U324 ( .A(n380), .B(n381), .Y(n382) );
  NAND2X2 U325 ( .A(n382), .B(n185), .Y(n183) );
  INVX2 U326 ( .A(n184), .Y(n380) );
  INVX2 U327 ( .A(n188), .Y(n381) );
  NOR2X2 U328 ( .A(A[13]), .B(B[13]), .Y(n184) );
  NAND2XL U329 ( .A(A[12]), .B(B[12]), .Y(n188) );
  NAND2X2 U330 ( .A(n383), .B(n384), .Y(n385) );
  NAND2X4 U331 ( .A(n385), .B(n124), .Y(n118) );
  INVXL U332 ( .A(n123), .Y(n383) );
  INVX2 U333 ( .A(n129), .Y(n384) );
  INVX2 U334 ( .A(n118), .Y(n120) );
  NAND2X4 U335 ( .A(n386), .B(n387), .Y(n388) );
  NAND2X4 U336 ( .A(n388), .B(n104), .Y(n102) );
  INVX2 U337 ( .A(n131), .Y(n386) );
  CLKINVX2 U338 ( .A(n103), .Y(n387) );
  AOI21X2 U339 ( .A0(n132), .A1(n168), .B0(n133), .Y(n131) );
  NAND2X1 U340 ( .A(n105), .B(n117), .Y(n103) );
  AOI21X2 U341 ( .A0(n105), .A1(n118), .B0(n106), .Y(n104) );
  INVX8 U342 ( .A(n102), .Y(n101) );
  INVX2 U343 ( .A(n96), .Y(n247) );
  AOI21X2 U344 ( .A0(n190), .A1(n182), .B0(n183), .Y(n181) );
  NOR2X2 U345 ( .A(A[21]), .B(B[21]), .Y(n123) );
  XOR2X4 U346 ( .A(n109), .B(n10), .Y(SUM[23]) );
  NAND2XL U347 ( .A(A[1]), .B(B[1]), .Y(n238) );
  OAI21X2 U348 ( .A0(n215), .A1(n213), .B0(n214), .Y(n212) );
  XNOR2X1 U349 ( .A(n149), .B(n15), .Y(SUM[18]) );
  CLKINVXL U350 ( .A(n123), .Y(n251) );
  NOR2X1 U351 ( .A(A[16]), .B(B[16]), .Y(n161) );
  NAND2X1 U352 ( .A(A[18]), .B(B[18]), .Y(n148) );
  OAI21X2 U353 ( .A0(n96), .A1(n100), .B0(n97), .Y(n91) );
  NOR2X1 U354 ( .A(n85), .B(n78), .Y(n76) );
  NAND2X1 U355 ( .A(n90), .B(n76), .Y(n70) );
  NOR2X1 U356 ( .A(n107), .B(n112), .Y(n105) );
  NAND2XL U357 ( .A(n54), .B(n38), .Y(n36) );
  AOI21X1 U358 ( .A0(n236), .A1(n411), .B0(n233), .Y(n231) );
  OAI21X1 U359 ( .A0(n223), .A1(n221), .B0(n222), .Y(n220) );
  XOR2X1 U360 ( .A(n197), .B(n22), .Y(SUM[11]) );
  OAI21X1 U361 ( .A0(n237), .A1(n240), .B0(n238), .Y(n236) );
  AOI21X2 U362 ( .A0(n204), .A1(n212), .B0(n205), .Y(n203) );
  OR2X1 U363 ( .A(A[11]), .B(B[11]), .Y(n408) );
  OR2X1 U364 ( .A(A[10]), .B(B[10]), .Y(n409) );
  XOR2X1 U365 ( .A(n101), .B(n9), .Y(SUM[24]) );
  XOR2X1 U366 ( .A(n211), .B(n25), .Y(SUM[8]) );
  XNOR2X1 U367 ( .A(n160), .B(n16), .Y(SUM[17]) );
  OAI21X1 U368 ( .A0(n167), .A1(n161), .B0(n162), .Y(n160) );
  XOR2X1 U369 ( .A(n116), .B(n11), .Y(SUM[22]) );
  NAND2X1 U370 ( .A(n250), .B(n115), .Y(n11) );
  XNOR2X1 U371 ( .A(n69), .B(n401), .Y(SUM[28]) );
  OAI21X1 U372 ( .A0(n101), .A1(n70), .B0(n71), .Y(n69) );
  XNOR2X1 U373 ( .A(n80), .B(n400), .Y(SUM[27]) );
  INVX2 U374 ( .A(n78), .Y(n245) );
  NAND2X1 U375 ( .A(A[17]), .B(B[17]), .Y(n159) );
  XNOR2X1 U376 ( .A(n51), .B(n3), .Y(SUM[30]) );
  INVX2 U377 ( .A(n70), .Y(n72) );
  NAND2X1 U378 ( .A(n256), .B(n390), .Y(n150) );
  OAI21X2 U379 ( .A0(n181), .A1(n169), .B0(n170), .Y(n168) );
  NAND2X1 U380 ( .A(n406), .B(n407), .Y(n169) );
  INVX2 U381 ( .A(n147), .Y(n254) );
  NOR2X1 U382 ( .A(A[18]), .B(B[18]), .Y(n147) );
  INVX2 U383 ( .A(n162), .Y(n164) );
  NOR2X1 U384 ( .A(A[20]), .B(B[20]), .Y(n128) );
  NAND2X1 U385 ( .A(A[20]), .B(B[20]), .Y(n129) );
  NAND2X1 U386 ( .A(A[22]), .B(B[22]), .Y(n115) );
  NOR2X2 U387 ( .A(A[25]), .B(B[25]), .Y(n96) );
  NAND2X1 U388 ( .A(A[25]), .B(B[25]), .Y(n97) );
  NOR2X1 U389 ( .A(A[26]), .B(B[26]), .Y(n85) );
  NOR2X1 U390 ( .A(n128), .B(n123), .Y(n117) );
  NOR2X1 U391 ( .A(A[22]), .B(B[22]), .Y(n112) );
  NOR2X1 U392 ( .A(A[23]), .B(B[23]), .Y(n107) );
  NAND2X1 U393 ( .A(A[26]), .B(B[26]), .Y(n86) );
  NOR2X1 U394 ( .A(A[27]), .B(B[27]), .Y(n78) );
  NOR2X1 U395 ( .A(n70), .B(n36), .Y(n399) );
  AND2X1 U396 ( .A(n403), .B(n240), .Y(SUM[0]) );
  OR2X1 U397 ( .A(A[4]), .B(B[4]), .Y(n391) );
  NAND2X1 U398 ( .A(A[16]), .B(B[16]), .Y(n162) );
  AOI21X2 U399 ( .A0(n130), .A1(n110), .B0(n111), .Y(n109) );
  OAI21X1 U400 ( .A0(n120), .A1(n112), .B0(n115), .Y(n111) );
  NAND2X1 U401 ( .A(n408), .B(n199), .Y(n392) );
  AND2X4 U402 ( .A(n392), .B(n196), .Y(n192) );
  NOR2X2 U403 ( .A(A[9]), .B(B[9]), .Y(n206) );
  CLKINVX2 U404 ( .A(n90), .Y(n88) );
  CLKINVX2 U405 ( .A(n190), .Y(n189) );
  NAND2XL U406 ( .A(n245), .B(n79), .Y(n400) );
  NAND2XL U407 ( .A(n83), .B(n86), .Y(n7) );
  XNOR2X1 U408 ( .A(n31), .B(n236), .Y(SUM[2]) );
  CLKINVX2 U409 ( .A(n219), .Y(n217) );
  NAND2X1 U410 ( .A(A[21]), .B(B[21]), .Y(n124) );
  NOR2X1 U411 ( .A(A[3]), .B(B[3]), .Y(n229) );
  CLKINVXL U412 ( .A(n68), .Y(n66) );
  NAND2X1 U413 ( .A(A[10]), .B(B[10]), .Y(n201) );
  NAND2X1 U414 ( .A(n243), .B(n61), .Y(n4) );
  NAND2XL U415 ( .A(n65), .B(n68), .Y(n401) );
  NAND2XL U416 ( .A(A[23]), .B(B[23]), .Y(n108) );
  CLKINVXL U417 ( .A(n213), .Y(n265) );
  XOR2XL U418 ( .A(n26), .B(n215), .Y(SUM[7]) );
  OAI21XL U419 ( .A0(n60), .A1(n68), .B0(n61), .Y(n55) );
  NOR2X1 U420 ( .A(n47), .B(n40), .Y(n38) );
  INVX3 U421 ( .A(n168), .Y(n167) );
  NAND2XL U422 ( .A(n406), .B(n174), .Y(n393) );
  INVX1 U423 ( .A(n174), .Y(n172) );
  INVX2 U424 ( .A(n161), .Y(n256) );
  CLKINVXL U425 ( .A(n91), .Y(n89) );
  AOI21X1 U426 ( .A0(n202), .A1(n409), .B0(n199), .Y(n197) );
  NAND2XL U427 ( .A(n90), .B(n83), .Y(n81) );
  NAND2XL U428 ( .A(n72), .B(n54), .Y(n52) );
  INVX2 U429 ( .A(n35), .Y(n398) );
  INVX2 U430 ( .A(n397), .Y(SUM[33]) );
  CLKINVXL U431 ( .A(n60), .Y(n243) );
  CLKINVXL U432 ( .A(n221), .Y(n267) );
  INVX2 U433 ( .A(n67), .Y(n65) );
  CLKINVXL U434 ( .A(n85), .Y(n83) );
  NAND2X1 U435 ( .A(A[7]), .B(B[7]), .Y(n214) );
  NAND2X1 U436 ( .A(A[27]), .B(B[27]), .Y(n79) );
  CLKINVXL U437 ( .A(n150), .Y(n152) );
  NAND2X1 U438 ( .A(n254), .B(n405), .Y(n134) );
  XNOR2X1 U439 ( .A(n140), .B(n14), .Y(SUM[19]) );
  NAND2XL U440 ( .A(n405), .B(n139), .Y(n14) );
  OAI21XL U441 ( .A0(n167), .A1(n150), .B0(n151), .Y(n149) );
  INVX1 U442 ( .A(n139), .Y(n137) );
  XOR2X1 U443 ( .A(n189), .B(n21), .Y(SUM[12]) );
  NAND2XL U444 ( .A(n260), .B(n188), .Y(n21) );
  CLKINVXL U445 ( .A(n187), .Y(n260) );
  NAND2BX1 U446 ( .AN(n107), .B(n108), .Y(n10) );
  NAND2X4 U447 ( .A(n251), .B(n124), .Y(n394) );
  CLKINVXL U448 ( .A(n99), .Y(n248) );
  OR2X4 U449 ( .A(A[15]), .B(B[15]), .Y(n406) );
  XNOR2X4 U450 ( .A(n98), .B(n395), .Y(SUM[25]) );
  NAND2X4 U451 ( .A(n247), .B(n97), .Y(n395) );
  NAND2XL U452 ( .A(A[15]), .B(B[15]), .Y(n174) );
  NAND2XL U453 ( .A(n408), .B(n196), .Y(n22) );
  XNOR2X1 U454 ( .A(n202), .B(n396), .Y(SUM[10]) );
  NAND2X1 U455 ( .A(n409), .B(n201), .Y(n396) );
  NAND2BXL U456 ( .AN(n209), .B(n210), .Y(n25) );
  NAND2BX1 U457 ( .AN(n40), .B(n41), .Y(n2) );
  CLKINVXL U458 ( .A(n212), .Y(n211) );
  NAND2XL U459 ( .A(n263), .B(n207), .Y(n24) );
  OAI21XL U460 ( .A0(n211), .A1(n209), .B0(n210), .Y(n208) );
  CLKINVXL U461 ( .A(n206), .Y(n263) );
  OAI2BB1X1 U462 ( .A0N(n399), .A1N(n102), .B0(n398), .Y(n397) );
  NAND2XL U463 ( .A(A[13]), .B(B[13]), .Y(n185) );
  INVXL U464 ( .A(n47), .Y(n242) );
  NOR2X2 U465 ( .A(n67), .B(n60), .Y(n54) );
  OAI21XL U466 ( .A0(n57), .A1(n47), .B0(n50), .Y(n46) );
  XNOR2XL U467 ( .A(n29), .B(n228), .Y(SUM[4]) );
  XOR2XL U468 ( .A(n402), .B(n220), .Y(SUM[6]) );
  AND2X1 U469 ( .A(n410), .B(n219), .Y(n402) );
  OAI21XL U470 ( .A0(n50), .A1(n40), .B0(n41), .Y(n39) );
  NOR2X2 U471 ( .A(A[7]), .B(B[7]), .Y(n213) );
  NAND2XL U472 ( .A(A[3]), .B(B[3]), .Y(n230) );
  NAND2XL U473 ( .A(A[4]), .B(B[4]), .Y(n227) );
  NAND2XL U474 ( .A(A[2]), .B(B[2]), .Y(n235) );
  OR2XL U475 ( .A(A[0]), .B(B[0]), .Y(n403) );
  INVX2 U476 ( .A(n397), .Y(SUM[34]) );
  INVX2 U477 ( .A(n397), .Y(SUM[35]) );
  INVX2 U478 ( .A(n397), .Y(SUM[32]) );
  NOR2X1 U479 ( .A(n150), .B(n134), .Y(n132) );
  INVX2 U480 ( .A(n179), .Y(n177) );
  INVX2 U481 ( .A(n148), .Y(n146) );
  NAND2XL U482 ( .A(n390), .B(n159), .Y(n16) );
  NAND2XL U483 ( .A(n152), .B(n254), .Y(n141) );
  XOR2X1 U484 ( .A(n167), .B(n17), .Y(SUM[16]) );
  NAND2XL U485 ( .A(n256), .B(n162), .Y(n17) );
  XOR2X1 U486 ( .A(n180), .B(n404), .Y(SUM[14]) );
  AND2X1 U487 ( .A(n407), .B(n179), .Y(n404) );
  NAND2XL U488 ( .A(n254), .B(n148), .Y(n15) );
  XNOR2X1 U489 ( .A(n130), .B(n13), .Y(SUM[20]) );
  NAND2X1 U490 ( .A(n252), .B(n129), .Y(n13) );
  CLKINVXL U491 ( .A(n128), .Y(n252) );
  INVX2 U492 ( .A(n129), .Y(n127) );
  OR2X1 U493 ( .A(A[19]), .B(B[19]), .Y(n405) );
  NOR2X2 U494 ( .A(n99), .B(n96), .Y(n90) );
  CLKINVXL U495 ( .A(n112), .Y(n250) );
  NAND2X1 U496 ( .A(A[19]), .B(B[19]), .Y(n139) );
  NAND2X1 U497 ( .A(A[14]), .B(B[14]), .Y(n179) );
  INVX2 U498 ( .A(n71), .Y(n73) );
  NAND2X1 U499 ( .A(n408), .B(n409), .Y(n191) );
  NOR2X1 U500 ( .A(n184), .B(n187), .Y(n182) );
  OR2X1 U501 ( .A(A[14]), .B(B[14]), .Y(n407) );
  NAND2X1 U502 ( .A(n248), .B(n100), .Y(n9) );
  NOR2X1 U503 ( .A(n206), .B(n209), .Y(n204) );
  OAI21X1 U504 ( .A0(n206), .A1(n210), .B0(n207), .Y(n205) );
  XNOR2X1 U505 ( .A(n208), .B(n24), .Y(SUM[9]) );
  NOR2BXL U506 ( .AN(n117), .B(n112), .Y(n110) );
  XNOR2X2 U507 ( .A(n186), .B(n20), .Y(SUM[13]) );
  NAND2X1 U508 ( .A(n259), .B(n185), .Y(n20) );
  OAI21X2 U509 ( .A0(n189), .A1(n187), .B0(n188), .Y(n186) );
  INVX2 U510 ( .A(n184), .Y(n259) );
  INVX2 U511 ( .A(n201), .Y(n199) );
  NOR2X1 U512 ( .A(n274), .B(n273), .Y(n40) );
  NOR2X1 U513 ( .A(A[24]), .B(B[24]), .Y(n99) );
  NAND2X1 U514 ( .A(A[24]), .B(B[24]), .Y(n100) );
  NAND2X1 U515 ( .A(n242), .B(n50), .Y(n3) );
  NOR2X1 U516 ( .A(A[12]), .B(B[12]), .Y(n187) );
  NOR2X1 U517 ( .A(A[8]), .B(B[8]), .Y(n209) );
  NAND2X1 U518 ( .A(A[11]), .B(B[11]), .Y(n196) );
  NAND2X1 U519 ( .A(A[9]), .B(B[9]), .Y(n207) );
  CLKINVXL U520 ( .A(n86), .Y(n84) );
  NAND2X1 U521 ( .A(A[8]), .B(B[8]), .Y(n210) );
  NOR2BXL U522 ( .AN(n54), .B(n47), .Y(n45) );
  AOI21X1 U523 ( .A0(n391), .A1(n228), .B0(n225), .Y(n223) );
  INVX2 U524 ( .A(n227), .Y(n225) );
  NAND2X1 U525 ( .A(n274), .B(n273), .Y(n41) );
  NAND2X1 U526 ( .A(n265), .B(n214), .Y(n26) );
  CLKINVXL U527 ( .A(n55), .Y(n57) );
  NAND2X1 U528 ( .A(n391), .B(n227), .Y(n29) );
  OAI21X1 U529 ( .A0(n231), .A1(n229), .B0(n230), .Y(n228) );
  XOR2X1 U530 ( .A(n28), .B(n223), .Y(SUM[5]) );
  NAND2X1 U531 ( .A(n267), .B(n222), .Y(n28) );
  XOR2X1 U532 ( .A(n30), .B(n231), .Y(SUM[3]) );
  NAND2X1 U533 ( .A(n269), .B(n230), .Y(n30) );
  INVX2 U534 ( .A(n229), .Y(n269) );
  NOR2X1 U535 ( .A(A[30]), .B(B[30]), .Y(n47) );
  INVX1 U536 ( .A(A[32]), .Y(n274) );
  INVX1 U537 ( .A(B[32]), .Y(n273) );
  NOR2X1 U538 ( .A(A[29]), .B(B[29]), .Y(n60) );
  NAND2X1 U539 ( .A(A[29]), .B(B[29]), .Y(n61) );
  OR2X1 U540 ( .A(A[6]), .B(B[6]), .Y(n410) );
  NAND2X1 U541 ( .A(A[30]), .B(B[30]), .Y(n50) );
  NOR2X1 U542 ( .A(A[28]), .B(B[28]), .Y(n67) );
  NAND2X1 U543 ( .A(A[6]), .B(B[6]), .Y(n219) );
  NAND2X1 U544 ( .A(A[28]), .B(B[28]), .Y(n68) );
  NOR2X1 U545 ( .A(A[5]), .B(B[5]), .Y(n221) );
  INVX2 U546 ( .A(n235), .Y(n233) );
  OR2X1 U547 ( .A(A[2]), .B(B[2]), .Y(n411) );
  NAND2X1 U548 ( .A(n411), .B(n235), .Y(n31) );
  NAND2X1 U549 ( .A(A[5]), .B(B[5]), .Y(n222) );
  NOR2X2 U550 ( .A(A[1]), .B(B[1]), .Y(n237) );
  XOR2X2 U551 ( .A(n32), .B(n240), .Y(SUM[1]) );
  NAND2X2 U552 ( .A(n271), .B(n238), .Y(n32) );
  INVX2 U553 ( .A(n237), .Y(n271) );
  NAND2X1 U554 ( .A(A[0]), .B(B[0]), .Y(n240) );
  OAI21X1 U555 ( .A0(n78), .A1(n86), .B0(n79), .Y(n77) );
  OAI21X1 U556 ( .A0(n107), .A1(n115), .B0(n108), .Y(n106) );
  OAI21X1 U557 ( .A0(n151), .A1(n134), .B0(n135), .Y(n133) );
  OAI21XL U558 ( .A0(n141), .A1(n167), .B0(n142), .Y(n140) );
  XNOR2X2 U559 ( .A(n42), .B(n2), .Y(SUM[31]) );
  NAND2X1 U560 ( .A(n45), .B(n72), .Y(n43) );
  AOI21XL U561 ( .A0(n73), .A1(n45), .B0(n46), .Y(n44) );
  OAI21XL U562 ( .A0(n43), .A1(n101), .B0(n44), .Y(n42) );
  OAI21X1 U563 ( .A0(n101), .A1(n52), .B0(n53), .Y(n51) );
  OAI21X1 U564 ( .A0(n101), .A1(n81), .B0(n82), .Y(n80) );
  OAI21X1 U565 ( .A0(n101), .A1(n63), .B0(n64), .Y(n62) );
  AOI21XL U566 ( .A0(n91), .A1(n83), .B0(n84), .Y(n82) );
  AOI21X2 U567 ( .A0(n76), .A1(n91), .B0(n77), .Y(n71) );
  AOI21X4 U568 ( .A0(n410), .A1(n220), .B0(n217), .Y(n215) );
  NAND2XL U569 ( .A(n72), .B(n65), .Y(n63) );
  OAI21X4 U570 ( .A0(n191), .A1(n203), .B0(n192), .Y(n190) );
  OAI21XL U571 ( .A0(n71), .A1(n36), .B0(n37), .Y(n35) );
endmodule


module PE_DW01_add_21 ( A, B, CI, SUM, CO );
  input [34:0] A;
  input [34:0] B;
  output [34:0] SUM;
  input CI;
  output CO;
  wire   n2, n5, n8, n9, n10, n12, n13, n15, n16, n17, n20, n21, n22, n24, n25,
         n26, n27, n28, n30, n31, n32, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n50, n51, n52, n53, n54, n55, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n115, n116, n117, n118, n120, n123, n124,
         n125, n127, n128, n129, n130, n131, n133, n134, n135, n137, n139,
         n140, n141, n142, n146, n148, n149, n150, n151, n152, n153, n157,
         n158, n159, n160, n161, n162, n164, n167, n168, n170, n172, n174,
         n175, n177, n179, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n194, n196, n197, n199, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n217, n219, n220, n221, n222, n223, n225, n227, n228, n229,
         n230, n231, n233, n235, n236, n237, n238, n240, n243, n245, n247,
         n248, n250, n251, n252, n255, n256, n259, n260, n263, n264, n265,
         n267, n273, n274, n379, n380, n381, n382, n383, n384, n385, n386,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414;

  AOI21X1 U7 ( .A0(n55), .A1(n38), .B0(n39), .Y(n37) );
  AOI21X1 U17 ( .A0(n73), .A1(n45), .B0(n46), .Y(n44) );
  NAND2X4 U56 ( .A(n90), .B(n76), .Y(n70) );
  OAI21X4 U75 ( .A0(n101), .A1(n88), .B0(n89), .Y(n87) );
  NOR2X2 U82 ( .A(n99), .B(n96), .Y(n90) );
  OAI21X4 U89 ( .A0(n101), .A1(n99), .B0(n100), .Y(n98) );
  OAI21X4 U96 ( .A0(n131), .A1(n103), .B0(n104), .Y(n102) );
  XOR2X4 U115 ( .A(n125), .B(n12), .Y(SUM[21]) );
  AOI21X1 U151 ( .A0(n153), .A1(n385), .B0(n146), .Y(n142) );
  AOI21X1 U239 ( .A0(n204), .A1(n212), .B0(n205), .Y(n203) );
  BUFX3 U311 ( .A(n109), .Y(n389) );
  AOI21X1 U312 ( .A0(n405), .A1(n146), .B0(n137), .Y(n135) );
  INVX1 U313 ( .A(n128), .Y(n252) );
  OR2X4 U314 ( .A(n150), .B(n134), .Y(n384) );
  NAND2X4 U315 ( .A(n379), .B(n380), .Y(n381) );
  NAND2X4 U316 ( .A(n381), .B(n124), .Y(n118) );
  INVX3 U317 ( .A(n123), .Y(n379) );
  INVX8 U318 ( .A(n129), .Y(n380) );
  NOR2X2 U319 ( .A(A[21]), .B(B[21]), .Y(n123) );
  NAND2X4 U320 ( .A(A[20]), .B(B[20]), .Y(n129) );
  NAND2XL U321 ( .A(A[21]), .B(B[21]), .Y(n124) );
  NAND2X1 U322 ( .A(n130), .B(n117), .Y(n382) );
  CLKINVXL U323 ( .A(n118), .Y(n383) );
  AND2X4 U324 ( .A(n382), .B(n383), .Y(n116) );
  NOR2X2 U325 ( .A(n128), .B(n123), .Y(n117) );
  XOR2X4 U326 ( .A(n116), .B(n393), .Y(SUM[22]) );
  NOR2X2 U327 ( .A(A[24]), .B(B[24]), .Y(n99) );
  AOI21X2 U328 ( .A0(n105), .A1(n118), .B0(n106), .Y(n104) );
  OAI21XL U329 ( .A0(n107), .A1(n115), .B0(n108), .Y(n106) );
  OAI21X4 U330 ( .A0(n96), .A1(n100), .B0(n97), .Y(n91) );
  NAND2X2 U331 ( .A(A[24]), .B(B[24]), .Y(n100) );
  NOR2X2 U332 ( .A(A[25]), .B(B[25]), .Y(n96) );
  OAI21X1 U333 ( .A0(n167), .A1(n161), .B0(n162), .Y(n160) );
  INVX3 U334 ( .A(n168), .Y(n167) );
  AOI21X1 U335 ( .A0(n413), .A1(n228), .B0(n225), .Y(n223) );
  NAND2X1 U336 ( .A(n251), .B(n124), .Y(n12) );
  NOR2X1 U337 ( .A(A[3]), .B(B[3]), .Y(n229) );
  AOI21X1 U338 ( .A0(n236), .A1(n414), .B0(n233), .Y(n231) );
  OAI21X1 U339 ( .A0(n215), .A1(n213), .B0(n214), .Y(n212) );
  OAI21X1 U340 ( .A0(n237), .A1(n240), .B0(n238), .Y(n236) );
  XOR2X1 U341 ( .A(n32), .B(n240), .Y(SUM[1]) );
  OAI21XL U342 ( .A0(n141), .A1(n167), .B0(n142), .Y(n140) );
  NAND2XL U343 ( .A(n152), .B(n385), .Y(n141) );
  XNOR2X1 U344 ( .A(n149), .B(n15), .Y(SUM[18]) );
  NOR2X1 U345 ( .A(A[16]), .B(B[16]), .Y(n161) );
  OR2X2 U346 ( .A(A[14]), .B(B[14]), .Y(n408) );
  NAND2XL U347 ( .A(A[14]), .B(B[14]), .Y(n179) );
  XNOR2X1 U348 ( .A(n42), .B(n2), .Y(SUM[31]) );
  OAI21X1 U349 ( .A0(n151), .A1(n134), .B0(n135), .Y(n133) );
  NOR2X2 U350 ( .A(A[1]), .B(B[1]), .Y(n237) );
  NAND2X1 U351 ( .A(A[1]), .B(B[1]), .Y(n238) );
  OAI21X1 U352 ( .A0(n231), .A1(n229), .B0(n230), .Y(n228) );
  XOR2X1 U353 ( .A(n30), .B(n231), .Y(SUM[3]) );
  AOI21X2 U354 ( .A0(n412), .A1(n220), .B0(n217), .Y(n215) );
  XOR2X1 U355 ( .A(n175), .B(n391), .Y(SUM[15]) );
  INVX2 U356 ( .A(n91), .Y(n89) );
  XOR2X1 U357 ( .A(n101), .B(n9), .Y(SUM[24]) );
  XNOR2X1 U358 ( .A(n31), .B(n236), .Y(SUM[2]) );
  NAND2X1 U359 ( .A(n414), .B(n235), .Y(n31) );
  XOR2X1 U360 ( .A(n211), .B(n25), .Y(SUM[8]) );
  NAND2X1 U361 ( .A(n250), .B(n115), .Y(n393) );
  INVX2 U362 ( .A(n112), .Y(n250) );
  XNOR2X2 U363 ( .A(n98), .B(n8), .Y(SUM[25]) );
  NAND2X1 U364 ( .A(n247), .B(n97), .Y(n8) );
  AOI21X1 U365 ( .A0(n73), .A1(n65), .B0(n66), .Y(n64) );
  NAND2X1 U366 ( .A(n72), .B(n65), .Y(n63) );
  XNOR2X1 U367 ( .A(n69), .B(n5), .Y(SUM[28]) );
  XNOR2X1 U368 ( .A(n80), .B(n398), .Y(SUM[27]) );
  OAI21X1 U369 ( .A0(n101), .A1(n81), .B0(n82), .Y(n80) );
  INVX2 U370 ( .A(n78), .Y(n245) );
  OAI21X1 U371 ( .A0(n191), .A1(n203), .B0(n192), .Y(n190) );
  NAND2X1 U372 ( .A(n410), .B(n411), .Y(n191) );
  INVX2 U373 ( .A(n161), .Y(n256) );
  NAND2X1 U374 ( .A(A[0]), .B(B[0]), .Y(n240) );
  XNOR2X1 U375 ( .A(n51), .B(n399), .Y(SUM[30]) );
  OAI21X1 U376 ( .A0(n101), .A1(n52), .B0(n53), .Y(n51) );
  XNOR2X1 U377 ( .A(n62), .B(n400), .Y(SUM[29]) );
  NAND2X1 U378 ( .A(n243), .B(n61), .Y(n400) );
  OAI21X1 U379 ( .A0(n101), .A1(n63), .B0(n64), .Y(n62) );
  INVX2 U380 ( .A(n60), .Y(n243) );
  INVX2 U381 ( .A(n71), .Y(n73) );
  NAND2X1 U382 ( .A(n256), .B(n255), .Y(n150) );
  OR2X1 U383 ( .A(A[18]), .B(B[18]), .Y(n385) );
  INVX2 U384 ( .A(n158), .Y(n255) );
  NOR2X1 U385 ( .A(A[17]), .B(B[17]), .Y(n158) );
  NAND2X1 U386 ( .A(A[16]), .B(B[16]), .Y(n162) );
  NAND2X1 U387 ( .A(A[17]), .B(B[17]), .Y(n159) );
  NAND2X1 U388 ( .A(n404), .B(n170), .Y(n168) );
  NAND2X1 U389 ( .A(n385), .B(n405), .Y(n134) );
  AOI21X2 U390 ( .A0(n255), .A1(n164), .B0(n157), .Y(n151) );
  INVX2 U391 ( .A(n159), .Y(n157) );
  INVX2 U392 ( .A(n162), .Y(n164) );
  NOR2X1 U393 ( .A(A[20]), .B(B[20]), .Y(n128) );
  NAND2X1 U394 ( .A(A[22]), .B(B[22]), .Y(n115) );
  NAND2X1 U395 ( .A(A[25]), .B(B[25]), .Y(n97) );
  NOR2X1 U396 ( .A(A[23]), .B(B[23]), .Y(n107) );
  NOR2X2 U397 ( .A(A[27]), .B(B[27]), .Y(n78) );
  NOR2X1 U398 ( .A(n70), .B(n36), .Y(n396) );
  XOR2X1 U399 ( .A(n197), .B(n22), .Y(SUM[11]) );
  AOI21X1 U400 ( .A0(n202), .A1(n411), .B0(n199), .Y(n197) );
  NAND2X1 U401 ( .A(n403), .B(n386), .Y(n404) );
  AOI21X1 U402 ( .A0(n403), .A1(n408), .B0(n177), .Y(n175) );
  AND2X1 U403 ( .A(n406), .B(n408), .Y(n386) );
  AOI21X1 U404 ( .A0(n190), .A1(n182), .B0(n183), .Y(n181) );
  NOR2X1 U405 ( .A(A[30]), .B(B[30]), .Y(n47) );
  AND2X1 U406 ( .A(n402), .B(n240), .Y(SUM[0]) );
  OAI21X1 U407 ( .A0(n223), .A1(n221), .B0(n222), .Y(n220) );
  INVX1 U408 ( .A(n221), .Y(n267) );
  NOR2X4 U409 ( .A(n384), .B(n167), .Y(n388) );
  NOR2X4 U410 ( .A(n388), .B(n133), .Y(n131) );
  AOI21X1 U411 ( .A0(n130), .A1(n110), .B0(n111), .Y(n109) );
  INVXL U412 ( .A(n99), .Y(n248) );
  NAND2XL U413 ( .A(n248), .B(n100), .Y(n9) );
  OAI21X1 U414 ( .A0(n101), .A1(n70), .B0(n71), .Y(n69) );
  AOI21X1 U415 ( .A0(n410), .A1(n199), .B0(n194), .Y(n192) );
  NAND2XL U416 ( .A(n245), .B(n79), .Y(n398) );
  OAI21XL U417 ( .A0(n167), .A1(n150), .B0(n151), .Y(n149) );
  NAND2XL U418 ( .A(A[27]), .B(B[27]), .Y(n79) );
  NAND2X2 U419 ( .A(n105), .B(n117), .Y(n103) );
  OR2X2 U420 ( .A(A[10]), .B(B[10]), .Y(n411) );
  NAND2XL U421 ( .A(A[10]), .B(B[10]), .Y(n201) );
  INVX4 U422 ( .A(n70), .Y(n72) );
  NAND2X1 U423 ( .A(A[18]), .B(B[18]), .Y(n148) );
  INVXL U424 ( .A(n67), .Y(n65) );
  OAI2BB1X1 U425 ( .A0N(n55), .A1N(n401), .B0(n50), .Y(n46) );
  NAND2XL U426 ( .A(n255), .B(n159), .Y(n16) );
  XNOR2X2 U427 ( .A(n160), .B(n16), .Y(SUM[17]) );
  AOI21X1 U428 ( .A0(n406), .A1(n177), .B0(n172), .Y(n170) );
  INVX2 U429 ( .A(n181), .Y(n403) );
  NAND2XL U430 ( .A(n256), .B(n162), .Y(n17) );
  NAND2X1 U431 ( .A(n252), .B(n129), .Y(n13) );
  AOI21X4 U432 ( .A0(n130), .A1(n252), .B0(n127), .Y(n125) );
  INVXL U433 ( .A(n123), .Y(n251) );
  INVX2 U434 ( .A(n35), .Y(n395) );
  INVX2 U435 ( .A(n394), .Y(SUM[33]) );
  INVX2 U436 ( .A(n219), .Y(n217) );
  INVX2 U437 ( .A(n227), .Y(n225) );
  NAND2XL U438 ( .A(n65), .B(n68), .Y(n5) );
  CLKINVXL U439 ( .A(n68), .Y(n66) );
  NAND2X1 U440 ( .A(n401), .B(n50), .Y(n399) );
  CLKINVXL U441 ( .A(n47), .Y(n401) );
  INVX2 U442 ( .A(n235), .Y(n233) );
  NAND2X1 U443 ( .A(A[3]), .B(B[3]), .Y(n230) );
  NAND2BXL U444 ( .AN(n237), .B(n238), .Y(n32) );
  XOR2X1 U445 ( .A(n167), .B(n17), .Y(SUM[16]) );
  XNOR2X2 U446 ( .A(n140), .B(n390), .Y(SUM[19]) );
  NAND2XL U447 ( .A(n405), .B(n139), .Y(n390) );
  CLKINVXL U448 ( .A(n190), .Y(n189) );
  NAND2XL U449 ( .A(n406), .B(n174), .Y(n391) );
  INVX1 U450 ( .A(n139), .Y(n137) );
  XOR2X1 U451 ( .A(n403), .B(n392), .Y(SUM[14]) );
  AND2X1 U452 ( .A(n408), .B(n179), .Y(n392) );
  CLKINVXL U453 ( .A(n129), .Y(n127) );
  NAND2BX1 U454 ( .AN(n107), .B(n108), .Y(n10) );
  XNOR2X1 U455 ( .A(n186), .B(n20), .Y(SUM[13]) );
  NAND2XL U456 ( .A(n259), .B(n185), .Y(n20) );
  OAI21XL U457 ( .A0(n189), .A1(n187), .B0(n188), .Y(n186) );
  CLKINVXL U458 ( .A(n184), .Y(n259) );
  NAND2XL U459 ( .A(n410), .B(n196), .Y(n22) );
  NAND2BX1 U460 ( .AN(n40), .B(n41), .Y(n2) );
  CLKINVXL U461 ( .A(n212), .Y(n211) );
  XOR2X1 U462 ( .A(n189), .B(n21), .Y(SUM[12]) );
  NAND2XL U463 ( .A(n260), .B(n188), .Y(n21) );
  CLKINVXL U464 ( .A(n187), .Y(n260) );
  XOR2X1 U465 ( .A(n202), .B(n407), .Y(SUM[10]) );
  OAI21XL U466 ( .A0(n211), .A1(n209), .B0(n210), .Y(n208) );
  CLKINVXL U467 ( .A(n206), .Y(n263) );
  OAI2BB1X1 U468 ( .A0N(n396), .A1N(n102), .B0(n395), .Y(n394) );
  NAND2XL U469 ( .A(A[11]), .B(B[11]), .Y(n196) );
  XNOR2X1 U470 ( .A(n397), .B(n228), .Y(SUM[4]) );
  NAND2XL U471 ( .A(n413), .B(n227), .Y(n397) );
  NAND2XL U472 ( .A(A[9]), .B(B[9]), .Y(n207) );
  XOR2XL U473 ( .A(n28), .B(n223), .Y(SUM[5]) );
  XOR2XL U474 ( .A(n26), .B(n215), .Y(SUM[7]) );
  NAND2XL U475 ( .A(n265), .B(n214), .Y(n26) );
  CLKINVXL U476 ( .A(n213), .Y(n265) );
  CLKINVXL U477 ( .A(n86), .Y(n84) );
  INVX1 U478 ( .A(n85), .Y(n83) );
  XNOR2XL U479 ( .A(n27), .B(n220), .Y(SUM[6]) );
  NAND2XL U480 ( .A(n412), .B(n219), .Y(n27) );
  OAI21XL U481 ( .A0(n60), .A1(n68), .B0(n61), .Y(n55) );
  NAND2BX1 U482 ( .AN(n229), .B(n230), .Y(n30) );
  NAND2XL U483 ( .A(A[30]), .B(B[30]), .Y(n50) );
  OR2XL U484 ( .A(A[0]), .B(B[0]), .Y(n402) );
  CLKINVXL U485 ( .A(n150), .Y(n152) );
  INVX2 U486 ( .A(n394), .Y(SUM[34]) );
  INVX2 U487 ( .A(n394), .Y(SUM[32]) );
  INVX2 U488 ( .A(n174), .Y(n172) );
  INVX2 U489 ( .A(n148), .Y(n146) );
  CLKINVXL U490 ( .A(n203), .Y(n202) );
  INVX2 U491 ( .A(n179), .Y(n177) );
  CLKINVXL U492 ( .A(n96), .Y(n247) );
  OAI21X1 U493 ( .A0(n184), .A1(n188), .B0(n185), .Y(n183) );
  NOR2X1 U494 ( .A(n184), .B(n187), .Y(n182) );
  OR2X1 U495 ( .A(A[19]), .B(B[19]), .Y(n405) );
  OR2X1 U496 ( .A(A[15]), .B(B[15]), .Y(n406) );
  INVX2 U497 ( .A(n196), .Y(n194) );
  AOI21X1 U498 ( .A0(n73), .A1(n54), .B0(n55), .Y(n53) );
  NAND2X1 U499 ( .A(A[19]), .B(B[19]), .Y(n139) );
  AND2X1 U500 ( .A(n411), .B(n201), .Y(n407) );
  NOR2BXL U501 ( .AN(n117), .B(n112), .Y(n110) );
  NAND2X1 U502 ( .A(A[15]), .B(B[15]), .Y(n174) );
  OAI21XL U503 ( .A0(n120), .A1(n112), .B0(n115), .Y(n111) );
  CLKINVXL U504 ( .A(n118), .Y(n120) );
  XNOR2X1 U505 ( .A(n208), .B(n24), .Y(SUM[9]) );
  NAND2X1 U506 ( .A(n263), .B(n207), .Y(n24) );
  NAND2X1 U507 ( .A(n264), .B(n210), .Y(n25) );
  INVX2 U508 ( .A(n209), .Y(n264) );
  OAI21XL U509 ( .A0(n43), .A1(n101), .B0(n44), .Y(n42) );
  INVX2 U510 ( .A(n201), .Y(n199) );
  NAND2XL U511 ( .A(n45), .B(n72), .Y(n43) );
  NOR2X1 U512 ( .A(n47), .B(n40), .Y(n38) );
  OAI21X1 U513 ( .A0(n50), .A1(n40), .B0(n41), .Y(n39) );
  NOR2X1 U514 ( .A(n67), .B(n60), .Y(n54) );
  NOR2X1 U515 ( .A(n274), .B(n273), .Y(n40) );
  XOR2X4 U516 ( .A(n87), .B(n409), .Y(SUM[26]) );
  AND2X1 U517 ( .A(n83), .B(n86), .Y(n409) );
  OAI21X2 U518 ( .A0(n78), .A1(n86), .B0(n79), .Y(n77) );
  NOR2X1 U519 ( .A(A[13]), .B(B[13]), .Y(n184) );
  NOR2X1 U520 ( .A(A[9]), .B(B[9]), .Y(n206) );
  OR2X4 U521 ( .A(A[11]), .B(B[11]), .Y(n410) );
  NOR2X1 U522 ( .A(A[12]), .B(B[12]), .Y(n187) );
  NAND2X1 U523 ( .A(A[8]), .B(B[8]), .Y(n210) );
  NOR2X1 U524 ( .A(A[8]), .B(B[8]), .Y(n209) );
  NAND2X1 U525 ( .A(A[13]), .B(B[13]), .Y(n185) );
  NAND2X1 U526 ( .A(A[23]), .B(B[23]), .Y(n108) );
  NAND2X1 U527 ( .A(n274), .B(n273), .Y(n41) );
  NAND2X1 U528 ( .A(n267), .B(n222), .Y(n28) );
  NAND2X1 U529 ( .A(A[12]), .B(B[12]), .Y(n188) );
  NOR2BXL U530 ( .AN(n54), .B(n47), .Y(n45) );
  NOR2X1 U531 ( .A(A[29]), .B(B[29]), .Y(n60) );
  INVX2 U532 ( .A(A[32]), .Y(n274) );
  NAND2X1 U533 ( .A(A[29]), .B(B[29]), .Y(n61) );
  NOR2X1 U534 ( .A(A[28]), .B(B[28]), .Y(n67) );
  INVX2 U535 ( .A(B[32]), .Y(n273) );
  NOR2X1 U536 ( .A(A[26]), .B(B[26]), .Y(n85) );
  OR2X1 U537 ( .A(A[6]), .B(B[6]), .Y(n412) );
  NOR2X1 U538 ( .A(A[5]), .B(B[5]), .Y(n221) );
  NAND2X1 U539 ( .A(A[26]), .B(B[26]), .Y(n86) );
  OR2X1 U540 ( .A(A[4]), .B(B[4]), .Y(n413) );
  NAND2X1 U541 ( .A(A[28]), .B(B[28]), .Y(n68) );
  NAND2X1 U542 ( .A(A[6]), .B(B[6]), .Y(n219) );
  NOR2X1 U543 ( .A(A[7]), .B(B[7]), .Y(n213) );
  NAND2X1 U544 ( .A(A[4]), .B(B[4]), .Y(n227) );
  OR2X1 U545 ( .A(A[2]), .B(B[2]), .Y(n414) );
  NAND2X1 U546 ( .A(A[7]), .B(B[7]), .Y(n214) );
  NAND2X1 U547 ( .A(A[2]), .B(B[2]), .Y(n235) );
  NAND2X1 U548 ( .A(A[5]), .B(B[5]), .Y(n222) );
  INVX2 U549 ( .A(n151), .Y(n153) );
  OAI21X1 U550 ( .A0(n206), .A1(n210), .B0(n207), .Y(n205) );
  NOR2X1 U551 ( .A(n206), .B(n209), .Y(n204) );
  XOR2X4 U552 ( .A(n389), .B(n10), .Y(SUM[23]) );
  INVX1 U553 ( .A(n90), .Y(n88) );
  NAND2X1 U554 ( .A(n90), .B(n83), .Y(n81) );
  NOR2X2 U555 ( .A(n107), .B(n112), .Y(n105) );
  OAI21XL U556 ( .A0(n71), .A1(n36), .B0(n37), .Y(n35) );
  AOI21XL U557 ( .A0(n91), .A1(n83), .B0(n84), .Y(n82) );
  XNOR2X1 U558 ( .A(n130), .B(n13), .Y(SUM[20]) );
  NAND2XL U559 ( .A(n385), .B(n148), .Y(n15) );
  INVX8 U560 ( .A(n102), .Y(n101) );
  NAND2XL U561 ( .A(n54), .B(n38), .Y(n36) );
  NAND2X1 U562 ( .A(n72), .B(n54), .Y(n52) );
  INVX4 U563 ( .A(n131), .Y(n130) );
  NOR2X4 U564 ( .A(n85), .B(n78), .Y(n76) );
  NOR2X4 U565 ( .A(A[22]), .B(B[22]), .Y(n112) );
  AOI21X4 U566 ( .A0(n76), .A1(n91), .B0(n77), .Y(n71) );
endmodule


module PE_DW01_add_22 ( A, B, CI, SUM, CO );
  input [37:0] A;
  input [37:0] B;
  output [37:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n6, n9, n12, n13, n14, n15, n16, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n33, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n57, n58, n59, n60, n62, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n98, n99, n100, n101, n102, n103, n104,
         n106, n110, n111, n112, n114, n116, n117, n118, n119, n120, n121,
         n122, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n141, n143, n144, n146, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n163, n165, n166, n168, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n198, n200, n201, n202, n203, n204, n206, n207, n208, n209, n210,
         n211, n212, n214, n216, n217, n219, n220, n221, n223, n229, n231,
         n232, n234, n237, n238, n241, n242, n245, n246, n248, n249, n250,
         n253, n254, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n385, n386, n387, n388, n389, n390, n391, n392, n393;

  XNOR2X4 U3 ( .A(n40), .B(n2), .Y(SUM[32]) );
  NAND2X4 U7 ( .A(n220), .B(n39), .Y(n2) );
  XNOR2X4 U71 ( .A(n91), .B(n9), .Y(SUM[25]) );
  NAND2X4 U106 ( .A(A[23]), .B(B[23]), .Y(n104) );
  XNOR2X4 U224 ( .A(n26), .B(n189), .Y(SUM[8]) );
  XOR2X4 U292 ( .A(n82), .B(n389), .Y(SUM[26]) );
  NOR2X4 U293 ( .A(A[21]), .B(B[21]), .Y(n120) );
  AOI21X2 U294 ( .A0(n78), .A1(n88), .B0(n79), .Y(n77) );
  NOR2X4 U295 ( .A(A[15]), .B(B[15]), .Y(n153) );
  OAI21X2 U296 ( .A0(n378), .A1(n83), .B0(n84), .Y(n82) );
  AOI21XL U297 ( .A0(n95), .A1(n87), .B0(n88), .Y(n84) );
  OR2X4 U298 ( .A(n43), .B(n41), .Y(n377) );
  INVX3 U299 ( .A(n44), .Y(n43) );
  NOR2X2 U300 ( .A(n92), .B(n76), .Y(n74) );
  INVX1 U301 ( .A(n172), .Y(n171) );
  INVX3 U302 ( .A(n73), .Y(n72) );
  OR2X4 U303 ( .A(A[22]), .B(B[22]), .Y(n369) );
  NAND2X1 U304 ( .A(A[20]), .B(B[20]), .Y(n126) );
  OR2X4 U305 ( .A(A[17]), .B(B[17]), .Y(n385) );
  AOI21X2 U306 ( .A0(n127), .A1(n232), .B0(n124), .Y(n122) );
  INVX4 U307 ( .A(n128), .Y(n127) );
  NAND2XL U308 ( .A(n110), .B(n94), .Y(n376) );
  NOR2X1 U309 ( .A(A[29]), .B(B[29]), .Y(n54) );
  AOI21XL U310 ( .A0(n44), .A1(n36), .B0(n37), .Y(SUM[34]) );
  NAND2XL U311 ( .A(n137), .B(n234), .Y(n375) );
  NAND2X4 U312 ( .A(n362), .B(n363), .Y(n364) );
  NAND2X4 U313 ( .A(n364), .B(n121), .Y(n119) );
  INVX2 U314 ( .A(n120), .Y(n362) );
  INVX2 U315 ( .A(n126), .Y(n363) );
  NAND2XL U316 ( .A(A[21]), .B(B[21]), .Y(n121) );
  AOI21X4 U317 ( .A0(n119), .A1(n369), .B0(n114), .Y(n112) );
  NAND2X1 U318 ( .A(n72), .B(n59), .Y(n365) );
  CLKINVXL U319 ( .A(n60), .Y(n366) );
  AND2X4 U320 ( .A(n365), .B(n366), .Y(n58) );
  NOR2X4 U321 ( .A(n70), .B(n65), .Y(n59) );
  XOR2X4 U322 ( .A(n58), .B(n383), .Y(SUM[29]) );
  NAND2X1 U323 ( .A(n72), .B(n68), .Y(n367) );
  INVX2 U324 ( .A(n69), .Y(n368) );
  AND2X4 U325 ( .A(n367), .B(n368), .Y(n67) );
  CLKINVXL U326 ( .A(n70), .Y(n68) );
  XOR2X4 U327 ( .A(n67), .B(n6), .Y(SUM[28]) );
  AOI21X2 U328 ( .A0(n385), .A1(n146), .B0(n141), .Y(n139) );
  XOR2X2 U329 ( .A(n51), .B(n4), .Y(SUM[30]) );
  AOI21X1 U330 ( .A0(n72), .A1(n52), .B0(n53), .Y(n51) );
  AOI21XL U331 ( .A0(n127), .A1(n118), .B0(n119), .Y(n117) );
  OAI21X1 U332 ( .A0(n131), .A1(n135), .B0(n132), .Y(n130) );
  NOR2X1 U333 ( .A(n131), .B(n134), .Y(n129) );
  OAI21X1 U334 ( .A0(n212), .A1(n210), .B0(n211), .Y(n209) );
  XNOR2X1 U335 ( .A(n33), .B(n217), .Y(SUM[1]) );
  NAND2X1 U336 ( .A(n223), .B(n57), .Y(n383) );
  CLKINVXL U337 ( .A(n54), .Y(n223) );
  NAND2X1 U338 ( .A(n221), .B(n42), .Y(n3) );
  CLKINVX2 U339 ( .A(n41), .Y(n221) );
  AOI21X1 U340 ( .A0(n173), .A1(n181), .B0(n174), .Y(n172) );
  NAND2XL U341 ( .A(A[1]), .B(B[1]), .Y(n216) );
  NAND2X1 U342 ( .A(n241), .B(n176), .Y(n23) );
  NAND2X1 U343 ( .A(A[18]), .B(B[18]), .Y(n135) );
  NOR2X1 U344 ( .A(A[20]), .B(B[20]), .Y(n125) );
  XNOR2X1 U345 ( .A(n31), .B(n209), .Y(SUM[3]) );
  INVXL U346 ( .A(n210), .Y(n250) );
  XOR2XL U347 ( .A(n25), .B(n184), .Y(SUM[9]) );
  AOI21XL U348 ( .A0(n149), .A1(n387), .B0(n146), .Y(n144) );
  NAND2X1 U349 ( .A(n229), .B(n104), .Y(n381) );
  AOI21X2 U350 ( .A0(n110), .A1(n74), .B0(n75), .Y(n73) );
  OAI21X1 U351 ( .A0(n204), .A1(n202), .B0(n203), .Y(n201) );
  OAI21X1 U352 ( .A0(n184), .A1(n182), .B0(n183), .Y(n181) );
  NOR2X2 U353 ( .A(A[11]), .B(B[11]), .Y(n175) );
  NAND2X1 U354 ( .A(A[3]), .B(B[3]), .Y(n208) );
  AOI21X2 U355 ( .A0(n209), .A1(n249), .B0(n206), .Y(n204) );
  INVX2 U356 ( .A(n208), .Y(n206) );
  INVX2 U357 ( .A(n100), .Y(n98) );
  NOR2X1 U358 ( .A(A[24]), .B(B[24]), .Y(n100) );
  INVX2 U359 ( .A(n216), .Y(n214) );
  NOR2X1 U360 ( .A(A[2]), .B(B[2]), .Y(n210) );
  NAND2X1 U361 ( .A(A[8]), .B(B[8]), .Y(n188) );
  NOR2X1 U362 ( .A(A[8]), .B(B[8]), .Y(n187) );
  INVX2 U363 ( .A(n192), .Y(n373) );
  XOR2X1 U364 ( .A(n27), .B(n192), .Y(SUM[7]) );
  AOI21X1 U365 ( .A0(n185), .A1(n193), .B0(n186), .Y(n184) );
  NOR2X1 U366 ( .A(n187), .B(n190), .Y(n185) );
  OAI21X1 U367 ( .A0(n187), .A1(n191), .B0(n188), .Y(n186) );
  XNOR2X1 U368 ( .A(n171), .B(n22), .Y(SUM[12]) );
  XOR2X1 U369 ( .A(n166), .B(n21), .Y(SUM[13]) );
  AND2X1 U370 ( .A(n372), .B(n170), .Y(n166) );
  XNOR2X1 U371 ( .A(n133), .B(n15), .Y(SUM[19]) );
  NAND2X1 U372 ( .A(n375), .B(n135), .Y(n133) );
  XNOR2X1 U373 ( .A(n127), .B(n14), .Y(SUM[20]) );
  OR2X1 U374 ( .A(A[16]), .B(B[16]), .Y(n387) );
  NOR2X1 U375 ( .A(n125), .B(n120), .Y(n118) );
  INVX2 U376 ( .A(n103), .Y(n229) );
  NOR2X2 U377 ( .A(A[28]), .B(B[28]), .Y(n65) );
  NAND2X1 U378 ( .A(n94), .B(n87), .Y(n83) );
  XOR2X1 U379 ( .A(n122), .B(n13), .Y(SUM[21]) );
  NAND2X1 U380 ( .A(n231), .B(n121), .Y(n13) );
  NOR2X1 U381 ( .A(A[30]), .B(B[30]), .Y(n49) );
  NOR2X1 U382 ( .A(n41), .B(n38), .Y(n36) );
  NAND2X1 U383 ( .A(n370), .B(n216), .Y(n33) );
  AOI21X1 U384 ( .A0(n370), .A1(n217), .B0(n214), .Y(n212) );
  AOI21X2 U385 ( .A0(n151), .A1(n159), .B0(n152), .Y(n150) );
  CLKINVXL U386 ( .A(n93), .Y(n95) );
  OAI21X2 U387 ( .A0(n150), .A1(n138), .B0(n139), .Y(n137) );
  INVX2 U388 ( .A(n110), .Y(n378) );
  OR2X1 U389 ( .A(A[1]), .B(B[1]), .Y(n370) );
  NAND2X1 U390 ( .A(n229), .B(n98), .Y(n92) );
  NOR2X1 U391 ( .A(A[18]), .B(B[18]), .Y(n134) );
  OR2X1 U392 ( .A(A[0]), .B(B[0]), .Y(n371) );
  XOR2X1 U393 ( .A(n43), .B(n3), .Y(SUM[31]) );
  NAND2X4 U394 ( .A(n377), .B(n42), .Y(n40) );
  NAND2X2 U395 ( .A(n376), .B(n93), .Y(n91) );
  INVX2 U396 ( .A(n159), .Y(n158) );
  NAND2X1 U397 ( .A(n388), .B(n390), .Y(n160) );
  AOI21X2 U398 ( .A0(n388), .A1(n168), .B0(n163), .Y(n161) );
  OAI21X2 U399 ( .A0(n153), .A1(n157), .B0(n154), .Y(n152) );
  NAND2XL U400 ( .A(n171), .B(n390), .Y(n372) );
  NOR2X2 U401 ( .A(n156), .B(n153), .Y(n151) );
  NAND2X2 U402 ( .A(n245), .B(n373), .Y(n374) );
  NAND2X2 U403 ( .A(n374), .B(n191), .Y(n189) );
  OAI21X4 U404 ( .A0(n128), .A1(n111), .B0(n112), .Y(n110) );
  OAI21X2 U405 ( .A0(n172), .A1(n160), .B0(n161), .Y(n159) );
  NAND2XL U406 ( .A(A[16]), .B(B[16]), .Y(n148) );
  INVX1 U407 ( .A(n165), .Y(n163) );
  NOR2X2 U408 ( .A(A[31]), .B(B[31]), .Y(n41) );
  INVX2 U409 ( .A(n181), .Y(n180) );
  INVX2 U410 ( .A(n125), .Y(n232) );
  NAND2X1 U411 ( .A(n254), .B(n253), .Y(n39) );
  NAND2BX1 U412 ( .AN(n65), .B(n66), .Y(n6) );
  NAND2X2 U413 ( .A(A[29]), .B(B[29]), .Y(n57) );
  XNOR2XL U414 ( .A(n392), .B(n212), .Y(SUM[2]) );
  AND2X1 U415 ( .A(n250), .B(n211), .Y(n392) );
  NAND2X4 U416 ( .A(A[31]), .B(B[31]), .Y(n42) );
  NAND2XL U417 ( .A(n385), .B(n143), .Y(n379) );
  XOR2X4 U418 ( .A(n378), .B(n381), .Y(SUM[23]) );
  NAND2XL U419 ( .A(n388), .B(n165), .Y(n21) );
  INVX4 U420 ( .A(n104), .Y(n106) );
  NOR2X1 U421 ( .A(n254), .B(n253), .Y(n38) );
  XNOR2X1 U422 ( .A(n72), .B(n382), .Y(SUM[27]) );
  NAND2XL U423 ( .A(n68), .B(n71), .Y(n382) );
  NAND2X1 U424 ( .A(A[2]), .B(B[2]), .Y(n211) );
  XOR2X1 U425 ( .A(n136), .B(n16), .Y(SUM[18]) );
  NAND2BX1 U426 ( .AN(n131), .B(n132), .Y(n15) );
  NAND2XL U427 ( .A(n232), .B(n126), .Y(n14) );
  XOR2X2 U428 ( .A(n144), .B(n379), .Y(SUM[17]) );
  XOR2X1 U429 ( .A(n149), .B(n380), .Y(SUM[16]) );
  AND2X1 U430 ( .A(n387), .B(n148), .Y(n380) );
  NAND2XL U431 ( .A(n237), .B(n154), .Y(n19) );
  CLKINVXL U432 ( .A(n153), .Y(n237) );
  XOR2X1 U433 ( .A(n158), .B(n20), .Y(SUM[14]) );
  NAND2XL U434 ( .A(n238), .B(n157), .Y(n20) );
  CLKINVXL U435 ( .A(n156), .Y(n238) );
  CLKINVXL U436 ( .A(n92), .Y(n94) );
  CLKINVXL U437 ( .A(n126), .Y(n124) );
  XOR2X1 U438 ( .A(n117), .B(n12), .Y(SUM[22]) );
  NAND2XL U439 ( .A(A[17]), .B(B[17]), .Y(n143) );
  INVX1 U440 ( .A(n170), .Y(n168) );
  CLKINVXL U441 ( .A(n175), .Y(n241) );
  NAND2XL U442 ( .A(n242), .B(n179), .Y(n24) );
  CLKINVXL U443 ( .A(n178), .Y(n242) );
  NAND2XL U444 ( .A(n390), .B(n170), .Y(n22) );
  NAND2BX1 U445 ( .AN(n182), .B(n183), .Y(n25) );
  OR2X4 U446 ( .A(A[13]), .B(B[13]), .Y(n388) );
  NAND2BX1 U447 ( .AN(n49), .B(n50), .Y(n4) );
  NAND2XL U448 ( .A(A[13]), .B(B[13]), .Y(n165) );
  NAND2XL U449 ( .A(A[22]), .B(B[22]), .Y(n116) );
  NAND2XL U450 ( .A(A[24]), .B(B[24]), .Y(n101) );
  OAI21X1 U451 ( .A0(n194), .A1(n196), .B0(n195), .Y(n193) );
  NAND2XL U452 ( .A(n245), .B(n191), .Y(n27) );
  CLKINVXL U453 ( .A(n190), .Y(n245) );
  NAND2BX1 U454 ( .AN(n187), .B(n188), .Y(n26) );
  CLKINVXL U455 ( .A(n60), .Y(n62) );
  XOR2XL U456 ( .A(n28), .B(n196), .Y(SUM[6]) );
  CLKINVXL U457 ( .A(n194), .Y(n246) );
  NAND2XL U458 ( .A(n248), .B(n203), .Y(n30) );
  CLKINVXL U459 ( .A(n202), .Y(n248) );
  XNOR2XL U460 ( .A(n29), .B(n201), .Y(SUM[5]) );
  NAND2XL U461 ( .A(A[9]), .B(B[9]), .Y(n183) );
  CLKINVXL U462 ( .A(n71), .Y(n69) );
  NAND2XL U463 ( .A(n249), .B(n208), .Y(n31) );
  NAND2X1 U464 ( .A(A[26]), .B(B[26]), .Y(n81) );
  OR2X2 U465 ( .A(A[5]), .B(B[5]), .Y(n391) );
  NAND2XL U466 ( .A(A[30]), .B(B[30]), .Y(n50) );
  NAND2XL U467 ( .A(A[5]), .B(B[5]), .Y(n200) );
  AND2X1 U468 ( .A(n371), .B(n219), .Y(SUM[0]) );
  CLKINVXL U469 ( .A(n150), .Y(n149) );
  CLKINVXL U470 ( .A(n137), .Y(n136) );
  INVX2 U471 ( .A(n393), .Y(SUM[37]) );
  INVX2 U472 ( .A(n393), .Y(SUM[36]) );
  INVX2 U473 ( .A(n393), .Y(SUM[35]) );
  INVX2 U474 ( .A(n393), .Y(SUM[33]) );
  NAND2X1 U475 ( .A(n385), .B(n387), .Y(n138) );
  INVX2 U476 ( .A(n143), .Y(n141) );
  INVX2 U477 ( .A(n148), .Y(n146) );
  XNOR2X1 U478 ( .A(n155), .B(n19), .Y(SUM[15]) );
  OAI21X1 U479 ( .A0(n158), .A1(n156), .B0(n157), .Y(n155) );
  NAND2XL U480 ( .A(n234), .B(n135), .Y(n16) );
  CLKINVXL U481 ( .A(n134), .Y(n234) );
  CLKINVXL U482 ( .A(SUM[34]), .Y(n393) );
  OAI21X1 U483 ( .A0(n42), .A1(n38), .B0(n39), .Y(n37) );
  CLKINVXL U484 ( .A(n38), .Y(n220) );
  INVX2 U485 ( .A(n116), .Y(n114) );
  INVX2 U486 ( .A(n101), .Y(n99) );
  INVX2 U487 ( .A(n90), .Y(n88) );
  NOR2X1 U488 ( .A(A[19]), .B(B[19]), .Y(n131) );
  CLKINVXL U489 ( .A(n120), .Y(n231) );
  XOR2X4 U490 ( .A(n102), .B(n386), .Y(SUM[24]) );
  AND2X1 U491 ( .A(n98), .B(n101), .Y(n386) );
  XNOR2X2 U492 ( .A(n177), .B(n23), .Y(SUM[11]) );
  NAND2X1 U493 ( .A(A[19]), .B(B[19]), .Y(n132) );
  NAND2X1 U494 ( .A(A[15]), .B(B[15]), .Y(n154) );
  NAND2XL U495 ( .A(n369), .B(n116), .Y(n12) );
  NOR2X1 U496 ( .A(A[14]), .B(B[14]), .Y(n156) );
  INVX2 U497 ( .A(n193), .Y(n192) );
  XOR2X1 U498 ( .A(n24), .B(n180), .Y(SUM[10]) );
  NAND2X1 U499 ( .A(A[14]), .B(B[14]), .Y(n157) );
  INVX2 U500 ( .A(A[33]), .Y(n254) );
  INVX2 U501 ( .A(B[33]), .Y(n253) );
  OAI21X2 U502 ( .A0(n65), .A1(n71), .B0(n66), .Y(n60) );
  INVX2 U503 ( .A(n81), .Y(n79) );
  NOR2BXL U504 ( .AN(n59), .B(n54), .Y(n52) );
  NAND2X2 U505 ( .A(A[25]), .B(B[25]), .Y(n90) );
  OAI21XL U506 ( .A0(n62), .A1(n54), .B0(n57), .Y(n53) );
  NOR2X1 U507 ( .A(A[10]), .B(B[10]), .Y(n178) );
  NOR2X1 U508 ( .A(A[9]), .B(B[9]), .Y(n182) );
  NAND2X2 U509 ( .A(A[11]), .B(B[11]), .Y(n176) );
  NAND2X1 U510 ( .A(A[10]), .B(B[10]), .Y(n179) );
  NAND2X1 U511 ( .A(n391), .B(n200), .Y(n29) );
  AOI21XL U512 ( .A0(n391), .A1(n201), .B0(n198), .Y(n196) );
  INVX2 U513 ( .A(n200), .Y(n198) );
  NAND2X1 U514 ( .A(n246), .B(n195), .Y(n28) );
  XOR2X2 U515 ( .A(n30), .B(n204), .Y(SUM[4]) );
  AND2X1 U516 ( .A(n78), .B(n81), .Y(n389) );
  OR2X1 U517 ( .A(A[12]), .B(B[12]), .Y(n390) );
  NAND2X1 U518 ( .A(A[12]), .B(B[12]), .Y(n170) );
  NOR2X1 U519 ( .A(A[27]), .B(B[27]), .Y(n70) );
  NAND2X1 U520 ( .A(A[27]), .B(B[27]), .Y(n71) );
  NAND2X1 U521 ( .A(A[28]), .B(B[28]), .Y(n66) );
  NOR2X1 U522 ( .A(A[4]), .B(B[4]), .Y(n202) );
  NOR2X1 U523 ( .A(A[6]), .B(B[6]), .Y(n194) );
  NAND2X1 U524 ( .A(A[7]), .B(B[7]), .Y(n191) );
  NOR2X1 U525 ( .A(A[7]), .B(B[7]), .Y(n190) );
  NAND2X1 U526 ( .A(A[6]), .B(B[6]), .Y(n195) );
  NAND2X1 U527 ( .A(A[4]), .B(B[4]), .Y(n203) );
  INVX2 U528 ( .A(n219), .Y(n217) );
  NAND2X1 U529 ( .A(A[0]), .B(B[0]), .Y(n219) );
  NAND2X2 U530 ( .A(n118), .B(n369), .Y(n111) );
  AOI21X1 U531 ( .A0(n47), .A1(n60), .B0(n48), .Y(n46) );
  OAI21X1 U532 ( .A0(n175), .A1(n179), .B0(n176), .Y(n174) );
  NOR2X1 U533 ( .A(n178), .B(n175), .Y(n173) );
  OAI21X4 U534 ( .A0(n378), .A1(n103), .B0(n104), .Y(n102) );
  NAND2XL U535 ( .A(n87), .B(n90), .Y(n9) );
  INVX4 U536 ( .A(n80), .Y(n78) );
  OAI21X2 U537 ( .A0(n73), .A1(n45), .B0(n46), .Y(n44) );
  NOR2X4 U538 ( .A(A[26]), .B(B[26]), .Y(n80) );
  OAI21X2 U539 ( .A0(n180), .A1(n178), .B0(n179), .Y(n177) );
  NAND2X1 U540 ( .A(n47), .B(n59), .Y(n45) );
  NOR2X2 U541 ( .A(n49), .B(n54), .Y(n47) );
  CLKINVX8 U542 ( .A(n89), .Y(n87) );
  NOR2X4 U543 ( .A(A[23]), .B(B[23]), .Y(n103) );
  NAND2X4 U544 ( .A(n87), .B(n78), .Y(n76) );
  NOR2X4 U545 ( .A(A[25]), .B(B[25]), .Y(n89) );
  OAI21XL U546 ( .A0(n49), .A1(n57), .B0(n50), .Y(n48) );
  NOR2X4 U547 ( .A(A[3]), .B(B[3]), .Y(n207) );
  OAI21X2 U548 ( .A0(n93), .A1(n76), .B0(n77), .Y(n75) );
  AOI21X4 U549 ( .A0(n98), .A1(n106), .B0(n99), .Y(n93) );
  AOI21X4 U550 ( .A0(n129), .A1(n137), .B0(n130), .Y(n128) );
  INVX4 U551 ( .A(n207), .Y(n249) );
endmodule


module PE_DW01_add_23 ( A, B, CI, SUM, CO );
  input [38:0] A;
  input [38:0] B;
  output [38:0] SUM;
  input CI;
  output CO;
  wire   n418, n3, n4, n5, n7, n8, n9, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n25, n26, n27, n28, n29, n30, n31, n33, n37, n38,
         n39, n40, n42, n44, n45, n46, n47, n50, n51, n52, n53, n54, n55, n56,
         n58, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n74,
         n75, n76, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n121, n123, n124, n125, n126, n127, n128, n129, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n148, n150, n151, n153, n155, n156, n157,
         n159, n161, n162, n163, n164, n165, n167, n168, n169, n170, n171,
         n172, n174, n176, n177, n179, n181, n182, n183, n185, n187, n188,
         n189, n190, n191, n193, n195, n196, n197, n198, n199, n201, n203,
         n204, n205, n206, n207, n209, n211, n212, n213, n214, n215, n217,
         n219, n220, n222, n225, n227, n228, n229, n231, n232, n233, n234,
         n236, n237, n238, n239, n243, n244, n248, n250, n252, n254, n257,
         n258, n369, n370, n371, n372, n373, n374, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n407;

  AOI21X1 U8 ( .A0(n376), .A1(n51), .B0(n42), .Y(n40) );
  XNOR2X4 U71 ( .A(n94), .B(n8), .Y(SUM[27]) );
  OAI21X4 U91 ( .A0(n100), .A1(n106), .B0(n101), .Y(n99) );
  NAND2X4 U103 ( .A(B[24]), .B(A[24]), .Y(n106) );
  AOI21X1 U139 ( .A0(n134), .A1(n237), .B0(n131), .Y(n129) );
  XOR2X4 U161 ( .A(n151), .B(n19), .Y(SUM[16]) );
  AOI21X1 U165 ( .A0(n392), .A1(n153), .B0(n148), .Y(n146) );
  OAI21X4 U190 ( .A0(n165), .A1(n163), .B0(n164), .Y(n162) );
  AOI21X1 U214 ( .A0(n397), .A1(n182), .B0(n179), .Y(n177) );
  XOR2X4 U258 ( .A(n31), .B(n207), .Y(SUM[4]) );
  NOR2X2 U276 ( .A(A[2]), .B(B[2]), .Y(n213) );
  NOR2X2 U297 ( .A(n127), .B(n132), .Y(n125) );
  OAI21X1 U298 ( .A0(n380), .A1(n96), .B0(n93), .Y(n91) );
  NAND2X2 U299 ( .A(A[32]), .B(B[32]), .Y(n53) );
  NAND2X2 U300 ( .A(B[19]), .B(A[19]), .Y(n133) );
  AOI21X1 U301 ( .A0(n90), .A1(n99), .B0(n91), .Y(n89) );
  NAND2X2 U302 ( .A(n90), .B(n98), .Y(n88) );
  NAND2X1 U303 ( .A(n371), .B(n56), .Y(n54) );
  OR2X4 U304 ( .A(B[21]), .B(A[21]), .Y(n377) );
  NAND2X2 U305 ( .A(n393), .B(n397), .Y(n171) );
  OAI21X2 U306 ( .A0(n143), .A1(n141), .B0(n142), .Y(n140) );
  NAND2X1 U307 ( .A(n392), .B(n150), .Y(n19) );
  OR2X4 U308 ( .A(B[16]), .B(A[16]), .Y(n392) );
  INVXL U309 ( .A(n117), .Y(n116) );
  NAND2X1 U310 ( .A(n125), .B(n377), .Y(n118) );
  OAI21X2 U311 ( .A0(n116), .A1(n114), .B0(n115), .Y(n113) );
  INVX1 U312 ( .A(n163), .Y(n243) );
  NAND2X4 U313 ( .A(B[28]), .B(A[28]), .Y(n85) );
  XOR2X2 U314 ( .A(n102), .B(n387), .Y(SUM[25]) );
  AOI21X2 U315 ( .A0(n107), .A1(n232), .B0(n104), .Y(n102) );
  NOR2X2 U316 ( .A(n95), .B(n380), .Y(n90) );
  OAI21X2 U317 ( .A0(n86), .A1(n66), .B0(n67), .Y(n65) );
  NAND2X2 U318 ( .A(n50), .B(n376), .Y(n39) );
  OR2X4 U319 ( .A(n257), .B(n258), .Y(n376) );
  CLKINVX4 U320 ( .A(n52), .Y(n50) );
  NOR2X2 U321 ( .A(A[32]), .B(B[32]), .Y(n52) );
  NAND2X1 U322 ( .A(A[31]), .B(B[31]), .Y(n64) );
  AOI21X2 U323 ( .A0(n393), .A1(n179), .B0(n174), .Y(n172) );
  INVX3 U324 ( .A(n108), .Y(n373) );
  NAND2X2 U325 ( .A(n369), .B(n370), .Y(n371) );
  INVX2 U326 ( .A(n86), .Y(n369) );
  INVXL U327 ( .A(n55), .Y(n370) );
  INVX4 U328 ( .A(n87), .Y(n86) );
  XNOR2X2 U329 ( .A(n54), .B(n3), .Y(SUM[32]) );
  NAND2X4 U330 ( .A(n372), .B(n373), .Y(n374) );
  NAND2X4 U331 ( .A(n374), .B(n89), .Y(n87) );
  CLKINVX3 U332 ( .A(n88), .Y(n372) );
  OAI2BB1X2 U333 ( .A0N(n87), .A1N(n75), .B0(n74), .Y(n72) );
  INVX2 U334 ( .A(n87), .Y(n385) );
  NOR2X2 U335 ( .A(B[27]), .B(A[27]), .Y(n380) );
  OAI21X4 U336 ( .A0(n63), .A1(n71), .B0(n64), .Y(n62) );
  OAI21X2 U337 ( .A0(n127), .A1(n133), .B0(n128), .Y(n126) );
  AOI21X2 U338 ( .A0(n117), .A1(n109), .B0(n110), .Y(n108) );
  OAI21X2 U339 ( .A0(n111), .A1(n115), .B0(n112), .Y(n110) );
  INVX1 U340 ( .A(B[34]), .Y(n257) );
  NAND2X1 U341 ( .A(A[1]), .B(B[1]), .Y(n219) );
  OAI21X1 U342 ( .A0(n215), .A1(n213), .B0(n214), .Y(n212) );
  AOI21X2 U343 ( .A0(n212), .A1(n378), .B0(n209), .Y(n207) );
  INVX2 U344 ( .A(n211), .Y(n209) );
  OAI21X1 U345 ( .A0(n145), .A1(n157), .B0(n146), .Y(n144) );
  NAND2XL U346 ( .A(n392), .B(n396), .Y(n145) );
  OAI21X1 U347 ( .A0(n207), .A1(n205), .B0(n206), .Y(n204) );
  NAND2X2 U348 ( .A(A[3]), .B(B[3]), .Y(n211) );
  NAND2X1 U349 ( .A(A[4]), .B(B[4]), .Y(n206) );
  NOR2X2 U350 ( .A(A[8]), .B(B[8]), .Y(n189) );
  INVX2 U351 ( .A(n183), .Y(n182) );
  NAND2X2 U352 ( .A(A[30]), .B(B[30]), .Y(n71) );
  OAI21X1 U353 ( .A0(n56), .A1(n39), .B0(n40), .Y(n38) );
  OAI21X2 U354 ( .A0(n118), .A1(n135), .B0(n119), .Y(n117) );
  AOI21X1 U355 ( .A0(n391), .A1(n220), .B0(n217), .Y(n215) );
  OAI21X2 U356 ( .A0(n191), .A1(n189), .B0(n190), .Y(n188) );
  AOI21X1 U357 ( .A0(n399), .A1(n204), .B0(n201), .Y(n199) );
  OR2X2 U358 ( .A(A[7]), .B(B[7]), .Y(n400) );
  OAI21X1 U359 ( .A0(n197), .A1(n199), .B0(n198), .Y(n196) );
  NOR2X1 U360 ( .A(A[12]), .B(B[12]), .Y(n168) );
  NAND2X1 U361 ( .A(B[13]), .B(A[13]), .Y(n164) );
  NOR2X2 U362 ( .A(B[13]), .B(A[13]), .Y(n163) );
  NOR2X1 U363 ( .A(B[19]), .B(A[19]), .Y(n132) );
  NOR2X1 U364 ( .A(B[20]), .B(A[20]), .Y(n127) );
  AOI21X2 U365 ( .A0(n136), .A1(n144), .B0(n137), .Y(n135) );
  OAI21X1 U366 ( .A0(n138), .A1(n142), .B0(n139), .Y(n137) );
  INVX2 U367 ( .A(n155), .Y(n153) );
  NAND2X1 U368 ( .A(n257), .B(n258), .Y(n44) );
  NAND2X1 U369 ( .A(n252), .B(n206), .Y(n31) );
  XNOR2X1 U370 ( .A(n25), .B(n182), .Y(SUM[10]) );
  NAND2X2 U371 ( .A(B[26]), .B(A[26]), .Y(n96) );
  NOR2X2 U372 ( .A(B[26]), .B(A[26]), .Y(n95) );
  XNOR2X1 U373 ( .A(n140), .B(n17), .Y(SUM[18]) );
  NAND2X1 U374 ( .A(B[21]), .B(A[21]), .Y(n123) );
  INVX2 U375 ( .A(n135), .Y(n134) );
  XNOR2X1 U376 ( .A(n65), .B(n4), .Y(SUM[31]) );
  XNOR2X1 U377 ( .A(n72), .B(n5), .Y(SUM[30]) );
  NAND2X1 U378 ( .A(n231), .B(n101), .Y(n387) );
  NAND2X1 U379 ( .A(n254), .B(n214), .Y(n33) );
  XNOR2X1 U380 ( .A(n26), .B(n188), .Y(SUM[9]) );
  BUFX2 U381 ( .A(SUM[38]), .Y(SUM[37]) );
  XNOR2X2 U382 ( .A(n113), .B(n12), .Y(SUM[23]) );
  AND2X1 U383 ( .A(n379), .B(n222), .Y(SUM[0]) );
  OR2X1 U384 ( .A(A[3]), .B(B[3]), .Y(n378) );
  XOR2X1 U385 ( .A(n33), .B(n215), .Y(SUM[2]) );
  OR2X1 U386 ( .A(A[0]), .B(B[0]), .Y(n379) );
  AOI21X1 U387 ( .A0(n37), .A1(n87), .B0(n38), .Y(n418) );
  OR2X2 U388 ( .A(B[9]), .B(A[9]), .Y(n395) );
  AOI21XL U389 ( .A0(n107), .A1(n98), .B0(n99), .Y(n97) );
  AOI21XL U390 ( .A0(n107), .A1(n98), .B0(n99), .Y(n381) );
  INVX2 U391 ( .A(n144), .Y(n143) );
  NAND2BX2 U392 ( .AN(n55), .B(n50), .Y(n46) );
  NAND2XL U393 ( .A(n75), .B(n68), .Y(n66) );
  INVX2 U394 ( .A(n157), .Y(n156) );
  AOI21X2 U395 ( .A0(n162), .A1(n398), .B0(n159), .Y(n157) );
  INVX1 U396 ( .A(n56), .Y(n58) );
  NOR2X2 U397 ( .A(B[29]), .B(A[29]), .Y(n81) );
  NOR2X2 U398 ( .A(n114), .B(n111), .Y(n109) );
  NAND2X1 U399 ( .A(A[12]), .B(B[12]), .Y(n169) );
  NOR2X1 U400 ( .A(n141), .B(n138), .Y(n136) );
  AOI21X2 U401 ( .A0(n126), .A1(n377), .B0(n121), .Y(n119) );
  INVX2 U402 ( .A(n108), .Y(n107) );
  NOR2X4 U403 ( .A(n382), .B(n168), .Y(n383) );
  NOR2X4 U404 ( .A(n383), .B(n167), .Y(n165) );
  CLKINVX4 U405 ( .A(n170), .Y(n382) );
  OAI21X2 U406 ( .A0(n171), .A1(n183), .B0(n172), .Y(n170) );
  INVX2 U407 ( .A(n168), .Y(n244) );
  INVX12 U408 ( .A(n169), .Y(n167) );
  NOR2X2 U409 ( .A(n70), .B(n63), .Y(n384) );
  NOR2X4 U410 ( .A(A[31]), .B(B[31]), .Y(n63) );
  AOI21X4 U411 ( .A0(n384), .A1(n76), .B0(n62), .Y(n56) );
  NOR2X1 U412 ( .A(n70), .B(n63), .Y(n61) );
  NOR2X2 U413 ( .A(B[28]), .B(A[28]), .Y(n84) );
  NOR2X1 U414 ( .A(n84), .B(n81), .Y(n75) );
  NOR2X4 U415 ( .A(B[24]), .B(A[24]), .Y(n105) );
  CLKINVX2 U416 ( .A(n44), .Y(n42) );
  CLKINVX2 U417 ( .A(n150), .Y(n148) );
  NAND2XL U418 ( .A(A[7]), .B(B[7]), .Y(n195) );
  OR2X1 U419 ( .A(A[1]), .B(B[1]), .Y(n391) );
  XOR2X1 U420 ( .A(n401), .B(n220), .Y(SUM[1]) );
  NAND2XL U421 ( .A(n236), .B(n128), .Y(n15) );
  INVX2 U422 ( .A(n123), .Y(n121) );
  XNOR2X1 U423 ( .A(n107), .B(n386), .Y(SUM[24]) );
  INVX2 U424 ( .A(n418), .Y(n407) );
  NOR2X1 U425 ( .A(n55), .B(n39), .Y(n37) );
  INVX4 U426 ( .A(n407), .Y(SUM[38]) );
  NAND2XL U427 ( .A(n393), .B(n176), .Y(n389) );
  OAI21X2 U428 ( .A0(n381), .A1(n95), .B0(n96), .Y(n94) );
  NAND2X2 U429 ( .A(B[25]), .B(A[25]), .Y(n101) );
  NAND2XL U430 ( .A(n225), .B(n64), .Y(n4) );
  XOR2X1 U431 ( .A(n83), .B(n394), .Y(SUM[29]) );
  NAND2XL U432 ( .A(n50), .B(n53), .Y(n3) );
  NAND2X1 U433 ( .A(A[8]), .B(B[8]), .Y(n190) );
  NAND2XL U434 ( .A(n237), .B(n133), .Y(n16) );
  NAND2XL U435 ( .A(n238), .B(n139), .Y(n17) );
  NAND2XL U436 ( .A(n239), .B(n142), .Y(n18) );
  CLKINVXL U437 ( .A(n141), .Y(n239) );
  CLKINVXL U438 ( .A(n138), .Y(n238) );
  NAND2XL U439 ( .A(B[20]), .B(A[20]), .Y(n128) );
  NAND2XL U440 ( .A(n232), .B(n106), .Y(n386) );
  XNOR2X2 U441 ( .A(n45), .B(n388), .Y(SUM[33]) );
  NAND2XL U442 ( .A(n376), .B(n44), .Y(n388) );
  NAND2XL U443 ( .A(n233), .B(n112), .Y(n12) );
  XOR2X1 U444 ( .A(n389), .B(n177), .Y(SUM[11]) );
  NAND2XL U445 ( .A(n398), .B(n161), .Y(n21) );
  NAND2XL U446 ( .A(n234), .B(n115), .Y(n13) );
  CLKINVXL U447 ( .A(n114), .Y(n234) );
  NAND2XL U448 ( .A(n395), .B(n187), .Y(n26) );
  NAND2BX1 U449 ( .AN(n95), .B(n96), .Y(n9) );
  OR2X4 U450 ( .A(B[11]), .B(A[11]), .Y(n393) );
  OR2X2 U451 ( .A(B[10]), .B(A[10]), .Y(n397) );
  NAND2XL U452 ( .A(B[14]), .B(A[14]), .Y(n161) );
  AOI21X1 U453 ( .A0(n58), .A1(n50), .B0(n51), .Y(n47) );
  NAND2XL U454 ( .A(B[11]), .B(A[11]), .Y(n176) );
  NAND2XL U455 ( .A(B[10]), .B(A[10]), .Y(n181) );
  NAND2X1 U456 ( .A(n248), .B(n190), .Y(n27) );
  NAND2XL U457 ( .A(n243), .B(n164), .Y(n22) );
  AND2X1 U458 ( .A(n227), .B(n82), .Y(n394) );
  NAND2X1 U459 ( .A(B[9]), .B(A[9]), .Y(n187) );
  CLKINVX2 U460 ( .A(n203), .Y(n201) );
  NAND2XL U461 ( .A(n250), .B(n198), .Y(n29) );
  CLKINVXL U462 ( .A(n197), .Y(n250) );
  CLKINVXL U463 ( .A(n380), .Y(n229) );
  CLKINVXL U464 ( .A(n70), .Y(n68) );
  NAND2XL U465 ( .A(n399), .B(n203), .Y(n30) );
  CLKINVXL U466 ( .A(n205), .Y(n252) );
  XOR2X1 U467 ( .A(n390), .B(n212), .Y(SUM[3]) );
  AND2X1 U468 ( .A(n378), .B(n211), .Y(n390) );
  AND2X1 U469 ( .A(n391), .B(n219), .Y(n401) );
  BUFX2 U470 ( .A(SUM[38]), .Y(SUM[34]) );
  XNOR2X1 U471 ( .A(n134), .B(n16), .Y(SUM[19]) );
  XOR2X1 U472 ( .A(n129), .B(n15), .Y(SUM[20]) );
  XOR2X1 U473 ( .A(n143), .B(n18), .Y(SUM[17]) );
  CLKINVXL U474 ( .A(n132), .Y(n237) );
  CLKINVXL U475 ( .A(n127), .Y(n236) );
  CLKINVXL U476 ( .A(n133), .Y(n131) );
  NAND2X1 U477 ( .A(n61), .B(n75), .Y(n55) );
  INVX2 U478 ( .A(n176), .Y(n174) );
  INVX2 U479 ( .A(n161), .Y(n159) );
  XNOR2X1 U480 ( .A(n156), .B(n20), .Y(SUM[15]) );
  NAND2X1 U481 ( .A(n396), .B(n155), .Y(n20) );
  NAND2X1 U482 ( .A(B[16]), .B(A[16]), .Y(n150) );
  XOR2X1 U483 ( .A(n124), .B(n14), .Y(SUM[21]) );
  NAND2XL U484 ( .A(n377), .B(n123), .Y(n14) );
  NOR2X1 U485 ( .A(B[17]), .B(A[17]), .Y(n141) );
  AOI21X2 U486 ( .A0(n395), .A1(n188), .B0(n185), .Y(n183) );
  INVX2 U487 ( .A(n187), .Y(n185) );
  NAND2X1 U488 ( .A(B[17]), .B(A[17]), .Y(n142) );
  NOR2X1 U489 ( .A(B[18]), .B(A[18]), .Y(n138) );
  NAND2X1 U490 ( .A(n397), .B(n181), .Y(n25) );
  INVX2 U491 ( .A(n181), .Y(n179) );
  CLKINVXL U492 ( .A(n111), .Y(n233) );
  NAND2X1 U493 ( .A(B[18]), .B(A[18]), .Y(n139) );
  INVX2 U494 ( .A(n105), .Y(n232) );
  CLKINVXL U495 ( .A(n100), .Y(n231) );
  CLKINVXL U496 ( .A(n106), .Y(n104) );
  XOR2X1 U497 ( .A(n116), .B(n13), .Y(SUM[22]) );
  INVX2 U498 ( .A(n53), .Y(n51) );
  NAND2X1 U499 ( .A(B[22]), .B(A[22]), .Y(n115) );
  NOR2X1 U500 ( .A(B[22]), .B(A[22]), .Y(n114) );
  XNOR2X1 U501 ( .A(n170), .B(n23), .Y(SUM[12]) );
  NAND2XL U502 ( .A(n244), .B(n169), .Y(n23) );
  XOR2XL U503 ( .A(n22), .B(n165), .Y(SUM[13]) );
  AOI21X2 U504 ( .A0(n400), .A1(n196), .B0(n193), .Y(n191) );
  INVX2 U505 ( .A(n195), .Y(n193) );
  XNOR2XL U506 ( .A(n30), .B(n204), .Y(SUM[5]) );
  XOR2XL U507 ( .A(n29), .B(n199), .Y(SUM[6]) );
  NAND2X1 U508 ( .A(B[23]), .B(A[23]), .Y(n112) );
  NAND2XL U509 ( .A(n68), .B(n71), .Y(n5) );
  CLKINVXL U510 ( .A(n71), .Y(n69) );
  XNOR2XL U511 ( .A(n28), .B(n196), .Y(SUM[7]) );
  NAND2X1 U512 ( .A(n400), .B(n195), .Y(n28) );
  NAND2X1 U513 ( .A(B[15]), .B(A[15]), .Y(n155) );
  OR2X4 U514 ( .A(B[15]), .B(A[15]), .Y(n396) );
  OR2X1 U515 ( .A(B[14]), .B(A[14]), .Y(n398) );
  XOR2XL U516 ( .A(n27), .B(n191), .Y(SUM[8]) );
  CLKINVXL U517 ( .A(n189), .Y(n248) );
  NOR2X2 U518 ( .A(B[30]), .B(A[30]), .Y(n70) );
  INVX2 U519 ( .A(A[34]), .Y(n258) );
  NAND2X1 U520 ( .A(B[29]), .B(A[29]), .Y(n82) );
  OR2X1 U521 ( .A(A[5]), .B(B[5]), .Y(n399) );
  NOR2X1 U522 ( .A(A[6]), .B(B[6]), .Y(n197) );
  NAND2X1 U523 ( .A(A[5]), .B(B[5]), .Y(n203) );
  INVX2 U524 ( .A(n222), .Y(n220) );
  NAND2X1 U525 ( .A(A[0]), .B(B[0]), .Y(n222) );
  BUFX2 U526 ( .A(SUM[38]), .Y(SUM[35]) );
  BUFX2 U527 ( .A(SUM[38]), .Y(SUM[36]) );
  NAND2X1 U528 ( .A(n229), .B(n93), .Y(n8) );
  CLKINVXL U529 ( .A(n81), .Y(n227) );
  INVX1 U530 ( .A(n84), .Y(n228) );
  INVXL U531 ( .A(n63), .Y(n225) );
  AOI21X1 U532 ( .A0(n76), .A1(n68), .B0(n69), .Y(n67) );
  INVX1 U533 ( .A(n76), .Y(n74) );
  NAND2X1 U534 ( .A(A[6]), .B(B[6]), .Y(n198) );
  XOR2X1 U535 ( .A(n97), .B(n9), .Y(SUM[26]) );
  AOI21XL U536 ( .A0(n134), .A1(n125), .B0(n126), .Y(n124) );
  OAI21X2 U537 ( .A0(n46), .A1(n86), .B0(n47), .Y(n45) );
  NAND2X1 U538 ( .A(B[27]), .B(A[27]), .Y(n93) );
  NAND2XL U539 ( .A(n228), .B(n85), .Y(n7) );
  NOR2X4 U540 ( .A(B[23]), .B(A[23]), .Y(n111) );
  XOR2X1 U541 ( .A(n385), .B(n7), .Y(SUM[28]) );
  OAI21X1 U542 ( .A0(n385), .A1(n84), .B0(n85), .Y(n83) );
  NOR2X4 U543 ( .A(n100), .B(n105), .Y(n98) );
  OAI21X4 U544 ( .A0(n81), .A1(n85), .B0(n82), .Y(n76) );
  AOI21X4 U545 ( .A0(n156), .A1(n396), .B0(n153), .Y(n151) );
  NOR2X4 U546 ( .A(B[25]), .B(A[25]), .Y(n100) );
  XNOR2XL U547 ( .A(n21), .B(n162), .Y(SUM[14]) );
  INVX2 U548 ( .A(n213), .Y(n254) );
  INVXL U549 ( .A(n219), .Y(n217) );
  NOR2X4 U550 ( .A(A[4]), .B(B[4]), .Y(n205) );
  NAND2X1 U551 ( .A(A[2]), .B(B[2]), .Y(n214) );
endmodule


module PE_DW01_add_17 ( A, B, CI, SUM, CO );
  input [33:0] A;
  input [33:0] B;
  output [33:0] SUM;
  input CI;
  output CO;
  wire   n1, n6, n7, n8, n9, n10, n11, n12, n13, n15, n16, n17, n18, n20, n21,
         n22, n25, n26, n27, n28, n29, n30, n31, n35, n36, n38, n40, n41, n43,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n64, n65, n66, n67, n68, n69, n71, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n129, n130, n131, n132, n134,
         n137, n138, n139, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n158, n160, n161,
         n162, n163, n164, n165, n166, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n185,
         n187, n188, n190, n192, n193, n194, n196, n198, n199, n200, n201,
         n202, n204, n206, n207, n208, n209, n210, n212, n214, n215, n216,
         n217, n218, n220, n222, n223, n224, n225, n227, n230, n231, n232,
         n234, n236, n238, n241, n242, n243, n245, n246, n247, n252, n254,
         n256, n258, n260, n261, n367, n368, n369, n370, n371, n372, n374,
         n375, n376, n377, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393;

  XOR2X4 U4 ( .A(n41), .B(n1), .Y(SUM[31]) );
  AOI21X1 U7 ( .A0(n389), .A1(n43), .B0(n38), .Y(n36) );
  XNOR2X4 U85 ( .A(n101), .B(n8), .Y(SUM[24]) );
  AOI21X1 U88 ( .A0(n105), .A1(n97), .B0(n98), .Y(n96) );
  OAI21X4 U96 ( .A0(n115), .A1(n102), .B0(n103), .Y(n101) );
  OAI21X4 U173 ( .A0(n155), .A1(n172), .B0(n156), .Y(n154) );
  AOI21XL U299 ( .A0(n144), .A1(n124), .B0(n125), .Y(n123) );
  NAND2X1 U300 ( .A(n86), .B(n79), .Y(n77) );
  NOR2X2 U301 ( .A(n151), .B(n148), .Y(n146) );
  OAI21X2 U302 ( .A0(n148), .A1(n152), .B0(n149), .Y(n147) );
  AOI21XL U303 ( .A0(n87), .A1(n79), .B0(n80), .Y(n78) );
  NAND2X1 U304 ( .A(n367), .B(n368), .Y(n369) );
  NAND2X2 U305 ( .A(n369), .B(n67), .Y(n65) );
  CLKINVXL U306 ( .A(n115), .Y(n367) );
  INVX1 U307 ( .A(n66), .Y(n368) );
  AOI21XL U308 ( .A0(n87), .A1(n68), .B0(n69), .Y(n67) );
  XOR2X4 U309 ( .A(n65), .B(n385), .Y(SUM[28]) );
  NAND2X4 U310 ( .A(n370), .B(n371), .Y(n372) );
  NAND2X2 U311 ( .A(n372), .B(n152), .Y(n150) );
  INVX3 U312 ( .A(n153), .Y(n370) );
  INVX12 U313 ( .A(n151), .Y(n371) );
  CLKINVX4 U314 ( .A(n154), .Y(n153) );
  XNOR2X2 U315 ( .A(n83), .B(n6), .Y(SUM[26]) );
  AOI21X2 U316 ( .A0(n90), .A1(n105), .B0(n91), .Y(n85) );
  OAI21X2 U317 ( .A0(n110), .A1(n114), .B0(n111), .Y(n105) );
  OAI21X2 U318 ( .A0(n115), .A1(n113), .B0(n114), .Y(n112) );
  XNOR2X2 U319 ( .A(n94), .B(n7), .Y(SUM[25]) );
  NAND2XL U320 ( .A(n234), .B(n93), .Y(n7) );
  AOI21X1 U321 ( .A0(n199), .A1(n387), .B0(n196), .Y(n194) );
  XOR2X1 U322 ( .A(n161), .B(n17), .Y(SUM[15]) );
  INVX2 U323 ( .A(n85), .Y(n87) );
  XOR2X1 U324 ( .A(n31), .B(n227), .Y(SUM[1]) );
  NAND2X1 U325 ( .A(n258), .B(n225), .Y(n31) );
  OR2X2 U326 ( .A(B[9]), .B(A[9]), .Y(n388) );
  XOR2X1 U327 ( .A(n139), .B(n13), .Y(SUM[19]) );
  CLKINVX2 U328 ( .A(n84), .Y(n86) );
  NOR2BX1 U329 ( .AN(n68), .B(n61), .Y(n59) );
  XOR2X1 U330 ( .A(n123), .B(n11), .Y(SUM[21]) );
  NAND2XL U331 ( .A(n238), .B(n122), .Y(n11) );
  AOI21XL U332 ( .A0(n87), .A1(n59), .B0(n60), .Y(n58) );
  OAI21XL U333 ( .A0(n71), .A1(n61), .B0(n64), .Y(n60) );
  INVXL U334 ( .A(n69), .Y(n71) );
  NOR2X1 U335 ( .A(n178), .B(n175), .Y(n173) );
  NAND2X1 U336 ( .A(B[26]), .B(A[26]), .Y(n82) );
  NOR2X1 U337 ( .A(B[1]), .B(A[1]), .Y(n224) );
  OR2X1 U338 ( .A(B[4]), .B(A[4]), .Y(n391) );
  XOR2X1 U339 ( .A(n180), .B(n21), .Y(SUM[11]) );
  OAI21X1 U340 ( .A0(n224), .A1(n227), .B0(n225), .Y(n223) );
  AOI21X1 U341 ( .A0(n392), .A1(n207), .B0(n204), .Y(n202) );
  XOR2X1 U342 ( .A(n130), .B(n12), .Y(SUM[20]) );
  NOR2X1 U343 ( .A(B[13]), .B(A[13]), .Y(n169) );
  NAND2X1 U344 ( .A(B[13]), .B(A[13]), .Y(n170) );
  NOR2X1 U345 ( .A(B[14]), .B(A[14]), .Y(n164) );
  OAI21X1 U346 ( .A0(n194), .A1(n182), .B0(n183), .Y(n181) );
  XOR2X2 U347 ( .A(n115), .B(n10), .Y(SUM[22]) );
  NAND2X1 U348 ( .A(n236), .B(n111), .Y(n9) );
  AND2X1 U349 ( .A(n231), .B(n64), .Y(n385) );
  XNOR2X1 U350 ( .A(n76), .B(n376), .Y(SUM[27]) );
  OAI21X1 U351 ( .A0(n115), .A1(n77), .B0(n78), .Y(n76) );
  XNOR2X1 U352 ( .A(n56), .B(n375), .Y(SUM[29]) );
  OAI21X1 U353 ( .A0(n115), .A1(n57), .B0(n58), .Y(n56) );
  INVX2 U354 ( .A(n54), .Y(n230) );
  AND2X1 U355 ( .A(n393), .B(n45), .Y(n384) );
  NOR2X1 U356 ( .A(B[23]), .B(A[23]), .Y(n110) );
  NAND2X1 U357 ( .A(B[23]), .B(A[23]), .Y(n111) );
  NAND2X1 U358 ( .A(B[20]), .B(A[20]), .Y(n129) );
  NOR2X1 U359 ( .A(n113), .B(n110), .Y(n104) );
  NOR2X1 U360 ( .A(B[28]), .B(A[28]), .Y(n61) );
  NOR2X1 U361 ( .A(B[29]), .B(A[29]), .Y(n54) );
  NAND2X1 U362 ( .A(B[28]), .B(A[28]), .Y(n64) );
  NAND2X1 U363 ( .A(B[29]), .B(A[29]), .Y(n55) );
  NOR2X1 U364 ( .A(n99), .B(n92), .Y(n90) );
  NOR2X1 U365 ( .A(B[25]), .B(A[25]), .Y(n92) );
  NAND2X1 U366 ( .A(B[25]), .B(A[25]), .Y(n93) );
  NOR2X1 U367 ( .A(B[26]), .B(A[26]), .Y(n81) );
  NOR2X2 U368 ( .A(B[20]), .B(A[20]), .Y(n126) );
  NOR2X2 U369 ( .A(B[21]), .B(A[21]), .Y(n121) );
  NAND2X1 U370 ( .A(n104), .B(n90), .Y(n84) );
  NOR2X1 U371 ( .A(n61), .B(n54), .Y(n52) );
  OAI21X1 U372 ( .A0(n92), .A1(n100), .B0(n93), .Y(n91) );
  AND2X1 U373 ( .A(n380), .B(n227), .Y(SUM[0]) );
  OAI21X2 U374 ( .A0(n115), .A1(n84), .B0(n85), .Y(n83) );
  XNOR2X2 U375 ( .A(n112), .B(n9), .Y(SUM[23]) );
  OAI21X2 U376 ( .A0(n115), .A1(n95), .B0(n96), .Y(n94) );
  INVX3 U377 ( .A(n145), .Y(n144) );
  NAND2BX1 U378 ( .AN(n178), .B(n179), .Y(n21) );
  OAI21X1 U379 ( .A0(n74), .A1(n82), .B0(n75), .Y(n69) );
  INVX2 U380 ( .A(n74), .Y(n232) );
  NOR2X1 U381 ( .A(n81), .B(n74), .Y(n68) );
  AOI21X2 U382 ( .A0(n173), .A1(n181), .B0(n174), .Y(n172) );
  AOI21X4 U383 ( .A0(n46), .A1(n393), .B0(n43), .Y(n41) );
  XOR2X1 U384 ( .A(n46), .B(n384), .Y(SUM[30]) );
  NAND2X1 U385 ( .A(B[24]), .B(A[24]), .Y(n100) );
  AOI21XL U386 ( .A0(n193), .A1(n388), .B0(n190), .Y(n188) );
  AOI21X1 U387 ( .A0(n386), .A1(n190), .B0(n185), .Y(n183) );
  NOR2X2 U388 ( .A(B[24]), .B(A[24]), .Y(n99) );
  NAND2XL U389 ( .A(B[4]), .B(A[4]), .Y(n214) );
  AOI21X1 U390 ( .A0(n52), .A1(n69), .B0(n53), .Y(n51) );
  INVX1 U391 ( .A(n187), .Y(n185) );
  NAND2XL U392 ( .A(n230), .B(n55), .Y(n375) );
  CLKINVXL U393 ( .A(n142), .Y(n241) );
  AOI21XL U394 ( .A0(n48), .A1(n116), .B0(n49), .Y(n47) );
  XOR2X1 U395 ( .A(n166), .B(n18), .Y(SUM[14]) );
  NAND2XL U396 ( .A(n242), .B(n149), .Y(n15) );
  CLKINVX2 U397 ( .A(n160), .Y(n158) );
  AOI21XL U398 ( .A0(n171), .A1(n246), .B0(n168), .Y(n166) );
  NAND2BXL U399 ( .AN(n113), .B(n114), .Y(n10) );
  INVX2 U400 ( .A(n36), .Y(n379) );
  NAND2BXL U401 ( .AN(n126), .B(n129), .Y(n12) );
  NAND2BX1 U402 ( .AN(n137), .B(n138), .Y(n13) );
  XOR2X1 U403 ( .A(n144), .B(n374), .Y(SUM[18]) );
  AND2X1 U404 ( .A(n241), .B(n143), .Y(n374) );
  CLKINVXL U405 ( .A(n151), .Y(n243) );
  OAI21XL U406 ( .A0(n134), .A1(n126), .B0(n129), .Y(n125) );
  CLKINVXL U407 ( .A(n143), .Y(n141) );
  NAND2X1 U408 ( .A(n59), .B(n86), .Y(n57) );
  NAND2X2 U409 ( .A(n381), .B(n162), .Y(n155) );
  NOR2X4 U410 ( .A(n126), .B(n121), .Y(n119) );
  OR2X4 U411 ( .A(B[15]), .B(A[15]), .Y(n381) );
  XOR2X1 U412 ( .A(n188), .B(n22), .Y(SUM[10]) );
  AOI21XL U413 ( .A0(n171), .A1(n162), .B0(n163), .Y(n161) );
  NAND2XL U414 ( .A(B[17]), .B(A[17]), .Y(n149) );
  NAND2XL U415 ( .A(B[15]), .B(A[15]), .Y(n160) );
  XOR2X1 U416 ( .A(n199), .B(n383), .Y(SUM[8]) );
  XOR2X1 U417 ( .A(n193), .B(n382), .Y(SUM[9]) );
  NAND2XL U418 ( .A(B[14]), .B(A[14]), .Y(n165) );
  OR2X4 U419 ( .A(B[10]), .B(A[10]), .Y(n386) );
  NAND2X1 U420 ( .A(n232), .B(n75), .Y(n376) );
  XOR2X1 U421 ( .A(n171), .B(n377), .Y(SUM[13]) );
  AND2X1 U422 ( .A(n246), .B(n170), .Y(n377) );
  CLKINVXL U423 ( .A(n169), .Y(n246) );
  XNOR2X1 U424 ( .A(n177), .B(n20), .Y(SUM[12]) );
  CLKINVXL U425 ( .A(n175), .Y(n247) );
  OR2X2 U426 ( .A(B[8]), .B(A[8]), .Y(n387) );
  NAND2XL U427 ( .A(B[10]), .B(A[10]), .Y(n187) );
  NAND2XL U428 ( .A(B[9]), .B(A[9]), .Y(n192) );
  NAND2XL U429 ( .A(B[8]), .B(A[8]), .Y(n198) );
  NAND2XL U430 ( .A(n392), .B(n206), .Y(n26) );
  CLKINVXL U431 ( .A(n216), .Y(n256) );
  XOR2XL U432 ( .A(n25), .B(n202), .Y(SUM[7]) );
  NAND2XL U433 ( .A(n252), .B(n201), .Y(n25) );
  CLKINVXL U434 ( .A(n200), .Y(n252) );
  AOI2BB1X1 U435 ( .A0N(n47), .A1N(n35), .B0(n379), .Y(SUM[33]) );
  XOR2XL U436 ( .A(n27), .B(n210), .Y(SUM[5]) );
  NAND2XL U437 ( .A(n254), .B(n209), .Y(n27) );
  CLKINVXL U438 ( .A(n208), .Y(n254) );
  NAND2XL U439 ( .A(B[12]), .B(A[12]), .Y(n176) );
  AOI21X1 U440 ( .A0(n223), .A1(n390), .B0(n220), .Y(n218) );
  INVX1 U441 ( .A(n222), .Y(n220) );
  NAND2XL U442 ( .A(B[30]), .B(A[30]), .Y(n45) );
  OR2XL U443 ( .A(B[0]), .B(A[0]), .Y(n380) );
  INVX2 U444 ( .A(n47), .Y(n46) );
  NOR2X1 U445 ( .A(n142), .B(n137), .Y(n131) );
  XNOR2X2 U446 ( .A(n150), .B(n15), .Y(SUM[17]) );
  OAI21X1 U447 ( .A0(n143), .A1(n137), .B0(n138), .Y(n132) );
  NAND2XL U448 ( .A(n104), .B(n97), .Y(n95) );
  CLKINVXL U449 ( .A(n194), .Y(n193) );
  CLKINVXL U450 ( .A(n104), .Y(n102) );
  NOR2BXL U451 ( .AN(n131), .B(n126), .Y(n124) );
  XOR2X1 U452 ( .A(n153), .B(n16), .Y(SUM[16]) );
  NAND2XL U453 ( .A(n243), .B(n152), .Y(n16) );
  CLKINVXL U454 ( .A(n132), .Y(n134) );
  AOI21X1 U455 ( .A0(n144), .A1(n241), .B0(n141), .Y(n139) );
  NAND2XL U456 ( .A(n86), .B(n68), .Y(n66) );
  CLKINVXL U457 ( .A(n92), .Y(n234) );
  CLKINVXL U458 ( .A(n110), .Y(n236) );
  NAND2X1 U459 ( .A(n97), .B(n100), .Y(n8) );
  CLKINVXL U460 ( .A(n105), .Y(n103) );
  NOR2X1 U461 ( .A(B[18]), .B(A[18]), .Y(n142) );
  INVX2 U462 ( .A(n100), .Y(n98) );
  NOR2X1 U463 ( .A(B[19]), .B(A[19]), .Y(n137) );
  NOR2X2 U464 ( .A(B[17]), .B(A[17]), .Y(n148) );
  INVX2 U465 ( .A(n99), .Y(n97) );
  NOR2X2 U466 ( .A(B[16]), .B(A[16]), .Y(n151) );
  NAND2X1 U467 ( .A(n386), .B(n388), .Y(n182) );
  NAND2X1 U468 ( .A(B[18]), .B(A[18]), .Y(n143) );
  NAND2XL U469 ( .A(n381), .B(n160), .Y(n17) );
  INVX2 U470 ( .A(n172), .Y(n171) );
  CLKINVXL U471 ( .A(n121), .Y(n238) );
  INVX2 U472 ( .A(n198), .Y(n196) );
  AND2X1 U473 ( .A(n388), .B(n192), .Y(n382) );
  AND2X1 U474 ( .A(n387), .B(n198), .Y(n383) );
  INVX2 U475 ( .A(n192), .Y(n190) );
  NAND2X1 U476 ( .A(n245), .B(n165), .Y(n18) );
  CLKINVXL U477 ( .A(n164), .Y(n245) );
  NAND2X1 U478 ( .A(B[19]), .B(A[19]), .Y(n138) );
  NAND2X1 U479 ( .A(n386), .B(n187), .Y(n22) );
  INVX2 U480 ( .A(n40), .Y(n38) );
  BUFX1 U481 ( .A(SUM[33]), .Y(SUM[32]) );
  NAND2XL U482 ( .A(n79), .B(n82), .Y(n6) );
  CLKINVXL U483 ( .A(n82), .Y(n80) );
  NAND2X1 U484 ( .A(B[21]), .B(A[21]), .Y(n122) );
  OAI21XL U485 ( .A0(n54), .A1(n64), .B0(n55), .Y(n53) );
  NAND2X1 U486 ( .A(B[22]), .B(A[22]), .Y(n114) );
  OAI21X1 U487 ( .A0(n175), .A1(n179), .B0(n176), .Y(n174) );
  OAI21X1 U488 ( .A0(n218), .A1(n216), .B0(n217), .Y(n215) );
  OAI21X1 U489 ( .A0(n210), .A1(n208), .B0(n209), .Y(n207) );
  AOI21X1 U490 ( .A0(n391), .A1(n215), .B0(n212), .Y(n210) );
  INVX2 U491 ( .A(n214), .Y(n212) );
  INVX2 U492 ( .A(n206), .Y(n204) );
  NOR2X2 U493 ( .A(n169), .B(n164), .Y(n162) );
  NOR2X1 U494 ( .A(B[22]), .B(A[22]), .Y(n113) );
  NAND2X1 U495 ( .A(n247), .B(n176), .Y(n20) );
  OAI21X1 U496 ( .A0(n180), .A1(n178), .B0(n179), .Y(n177) );
  NOR2X1 U497 ( .A(B[11]), .B(A[11]), .Y(n178) );
  NAND2X1 U498 ( .A(B[11]), .B(A[11]), .Y(n179) );
  XOR2X1 U499 ( .A(n29), .B(n218), .Y(SUM[3]) );
  NAND2X1 U500 ( .A(n256), .B(n217), .Y(n29) );
  NAND2X1 U501 ( .A(n389), .B(n40), .Y(n1) );
  XNOR2X1 U502 ( .A(n28), .B(n215), .Y(SUM[4]) );
  NAND2X1 U503 ( .A(n391), .B(n214), .Y(n28) );
  NAND2X1 U504 ( .A(n393), .B(n389), .Y(n35) );
  CLKINVXL U505 ( .A(n81), .Y(n79) );
  CLKINVXL U506 ( .A(n170), .Y(n168) );
  INVX2 U507 ( .A(n45), .Y(n43) );
  OR2X1 U508 ( .A(n261), .B(n260), .Y(n389) );
  NAND2X1 U509 ( .A(n261), .B(n260), .Y(n40) );
  NOR2X1 U510 ( .A(B[27]), .B(A[27]), .Y(n74) );
  NAND2X1 U511 ( .A(B[27]), .B(A[27]), .Y(n75) );
  NOR2X1 U512 ( .A(B[7]), .B(A[7]), .Y(n200) );
  NOR2X1 U513 ( .A(B[3]), .B(A[3]), .Y(n216) );
  XNOR2X1 U514 ( .A(n30), .B(n223), .Y(SUM[2]) );
  NAND2X1 U515 ( .A(n390), .B(n222), .Y(n30) );
  OR2X1 U516 ( .A(B[2]), .B(A[2]), .Y(n390) );
  OR2X1 U517 ( .A(B[6]), .B(A[6]), .Y(n392) );
  NOR2X1 U518 ( .A(B[5]), .B(A[5]), .Y(n208) );
  NOR2X1 U519 ( .A(B[12]), .B(A[12]), .Y(n175) );
  NAND2X1 U520 ( .A(B[2]), .B(A[2]), .Y(n222) );
  NAND2X1 U521 ( .A(B[6]), .B(A[6]), .Y(n206) );
  NAND2X1 U522 ( .A(B[3]), .B(A[3]), .Y(n217) );
  NAND2X1 U523 ( .A(B[5]), .B(A[5]), .Y(n209) );
  NAND2X1 U524 ( .A(B[7]), .B(A[7]), .Y(n201) );
  OR2X1 U525 ( .A(B[30]), .B(A[30]), .Y(n393) );
  INVX2 U526 ( .A(B[32]), .Y(n260) );
  INVX2 U527 ( .A(A[32]), .Y(n261) );
  NAND2X1 U528 ( .A(B[1]), .B(A[1]), .Y(n225) );
  NAND2X1 U529 ( .A(B[0]), .B(A[0]), .Y(n227) );
  AOI21XL U530 ( .A0(n144), .A1(n131), .B0(n132), .Y(n130) );
  INVX2 U531 ( .A(n181), .Y(n180) );
  INVX2 U532 ( .A(n148), .Y(n242) );
  OAI21X1 U533 ( .A0(n121), .A1(n129), .B0(n122), .Y(n120) );
  NAND2X2 U534 ( .A(B[16]), .B(A[16]), .Y(n152) );
  INVX2 U535 ( .A(n61), .Y(n231) );
  AOI21X1 U536 ( .A0(n119), .A1(n132), .B0(n120), .Y(n118) );
  NAND2X1 U537 ( .A(n119), .B(n131), .Y(n117) );
  OAI21X1 U538 ( .A0(n85), .A1(n50), .B0(n51), .Y(n49) );
  NAND2X1 U539 ( .A(n68), .B(n52), .Y(n50) );
  OAI21X2 U540 ( .A0(n164), .A1(n170), .B0(n165), .Y(n163) );
  OAI21X4 U541 ( .A0(n117), .A1(n145), .B0(n118), .Y(n116) );
  AOI21X2 U542 ( .A0(n381), .A1(n163), .B0(n158), .Y(n156) );
  XNOR2X1 U543 ( .A(n26), .B(n207), .Y(SUM[6]) );
  INVX8 U544 ( .A(n116), .Y(n115) );
  NOR2X1 U545 ( .A(n84), .B(n50), .Y(n48) );
  INVX2 U546 ( .A(n224), .Y(n258) );
  AOI21X4 U547 ( .A0(n146), .A1(n154), .B0(n147), .Y(n145) );
  OAI21X2 U548 ( .A0(n202), .A1(n200), .B0(n201), .Y(n199) );
endmodule


module PE_DW01_add_20 ( A, B, CI, SUM, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] SUM;
  input CI;
  output CO;
  wire   n2, n4, n5, n6, n7, n8, n9, n12, n15, n16, n17, n21, n25, n26, n27,
         n28, n29, n30, n31, n34, n35, n37, n39, n40, n41, n42, n43, n44, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n64, n65, n66, n67, n68, n69, n71, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n90, n91, n92, n93, n94, n96, n97,
         n98, n99, n100, n101, n103, n104, n105, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n129, n130, n131, n132, n133, n134, n137, n138, n139, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n158, n160, n161, n162, n163, n164, n165,
         n166, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n185, n187, n188, n190, n192,
         n193, n194, n196, n198, n199, n200, n201, n202, n204, n206, n207,
         n208, n209, n210, n212, n214, n215, n216, n217, n218, n220, n222,
         n223, n224, n225, n227, n230, n231, n234, n236, n237, n238, n239,
         n240, n241, n242, n243, n245, n246, n247, n248, n260, n261, n366,
         n367, n368, n370, n371, n372, n373, n374, n375, n376, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395;

  AOI21X1 U5 ( .A0(n390), .A1(n44), .B0(n37), .Y(n35) );
  NOR2X2 U28 ( .A(n61), .B(n54), .Y(n52) );
  XNOR2X4 U60 ( .A(n83), .B(n6), .Y(SUM[26]) );
  NOR2X2 U68 ( .A(B[26]), .B(A[26]), .Y(n81) );
  AOI21X1 U87 ( .A0(n105), .A1(n97), .B0(n98), .Y(n96) );
  NOR2X2 U102 ( .A(n113), .B(n110), .Y(n104) );
  AOI21X1 U182 ( .A0(n171), .A1(n162), .B0(n163), .Y(n161) );
  AOI21X1 U190 ( .A0(n171), .A1(n246), .B0(n168), .Y(n166) );
  AOI21X1 U224 ( .A0(n193), .A1(n389), .B0(n190), .Y(n188) );
  OAI21X1 U298 ( .A0(n194), .A1(n182), .B0(n183), .Y(n181) );
  INVX2 U299 ( .A(n85), .Y(n87) );
  XNOR2X2 U300 ( .A(n112), .B(n9), .Y(SUM[23]) );
  AOI21X2 U301 ( .A0(n119), .A1(n132), .B0(n120), .Y(n118) );
  OAI21X2 U302 ( .A0(n143), .A1(n137), .B0(n138), .Y(n132) );
  AOI21X1 U303 ( .A0(n144), .A1(n131), .B0(n132), .Y(n130) );
  NAND2XL U304 ( .A(n388), .B(n389), .Y(n182) );
  NAND2X4 U305 ( .A(n366), .B(n367), .Y(n368) );
  NAND2X4 U306 ( .A(n368), .B(n156), .Y(n154) );
  INVX4 U307 ( .A(n155), .Y(n366) );
  INVX2 U308 ( .A(n172), .Y(n367) );
  NAND2X2 U309 ( .A(n385), .B(n162), .Y(n155) );
  AOI21X2 U310 ( .A0(n385), .A1(n163), .B0(n158), .Y(n156) );
  OAI21X2 U311 ( .A0(n148), .A1(n152), .B0(n149), .Y(n147) );
  NOR2X2 U312 ( .A(B[17]), .B(A[17]), .Y(n148) );
  NOR2X2 U313 ( .A(B[16]), .B(A[16]), .Y(n151) );
  AOI21X2 U314 ( .A0(n90), .A1(n105), .B0(n91), .Y(n85) );
  NOR2X2 U315 ( .A(n99), .B(n92), .Y(n90) );
  NOR2X1 U316 ( .A(B[1]), .B(A[1]), .Y(n224) );
  XNOR2X1 U317 ( .A(n94), .B(n7), .Y(SUM[25]) );
  NAND2XL U318 ( .A(n234), .B(n93), .Y(n7) );
  AOI21X1 U319 ( .A0(n223), .A1(n391), .B0(n220), .Y(n218) );
  OR2X1 U320 ( .A(B[2]), .B(A[2]), .Y(n391) );
  XOR2X1 U321 ( .A(n31), .B(n227), .Y(SUM[1]) );
  XNOR2X1 U322 ( .A(n166), .B(n371), .Y(SUM[14]) );
  AND2X2 U323 ( .A(n245), .B(n165), .Y(n371) );
  NOR2BX1 U324 ( .AN(n68), .B(n61), .Y(n59) );
  INVX2 U325 ( .A(n84), .Y(n86) );
  XOR2X1 U326 ( .A(n123), .B(n373), .Y(SUM[21]) );
  CLKINVXL U327 ( .A(n121), .Y(n238) );
  NAND2X1 U328 ( .A(B[29]), .B(A[29]), .Y(n55) );
  NAND2X1 U329 ( .A(n104), .B(n90), .Y(n84) );
  XOR2X2 U330 ( .A(n47), .B(n2), .Y(SUM[30]) );
  OAI21XL U331 ( .A0(n47), .A1(n41), .B0(n42), .Y(n40) );
  AOI21X1 U332 ( .A0(n173), .A1(n181), .B0(n174), .Y(n172) );
  OAI21X1 U333 ( .A0(n175), .A1(n179), .B0(n176), .Y(n174) );
  NOR2X1 U334 ( .A(n178), .B(n175), .Y(n173) );
  OAI21X1 U335 ( .A0(n218), .A1(n216), .B0(n217), .Y(n215) );
  XOR2X1 U336 ( .A(n180), .B(n21), .Y(SUM[11]) );
  NOR2X1 U337 ( .A(B[12]), .B(A[12]), .Y(n175) );
  NOR2X1 U338 ( .A(B[11]), .B(A[11]), .Y(n178) );
  NAND2X1 U339 ( .A(B[11]), .B(A[11]), .Y(n179) );
  NOR2X1 U340 ( .A(n169), .B(n164), .Y(n162) );
  XOR2X1 U341 ( .A(n29), .B(n218), .Y(SUM[3]) );
  NOR2X1 U342 ( .A(B[7]), .B(A[7]), .Y(n200) );
  AOI21X1 U343 ( .A0(n392), .A1(n207), .B0(n204), .Y(n202) );
  OR2X1 U344 ( .A(B[8]), .B(A[8]), .Y(n387) );
  OAI21X1 U345 ( .A0(n202), .A1(n200), .B0(n201), .Y(n199) );
  XOR2X1 U346 ( .A(n130), .B(n12), .Y(SUM[20]) );
  NAND2X1 U347 ( .A(B[26]), .B(A[26]), .Y(n82) );
  NOR2X2 U348 ( .A(B[25]), .B(A[25]), .Y(n92) );
  NAND2X1 U349 ( .A(B[25]), .B(A[25]), .Y(n93) );
  XNOR2X1 U350 ( .A(n30), .B(n223), .Y(SUM[2]) );
  XNOR2X1 U351 ( .A(n65), .B(n4), .Y(SUM[28]) );
  XNOR2X1 U352 ( .A(n76), .B(n5), .Y(SUM[27]) );
  NAND2X1 U353 ( .A(n230), .B(n55), .Y(n379) );
  INVX2 U354 ( .A(n54), .Y(n230) );
  NOR2X1 U355 ( .A(n84), .B(n50), .Y(n48) );
  AND2X1 U356 ( .A(n381), .B(n227), .Y(SUM[0]) );
  OR2X1 U357 ( .A(B[4]), .B(A[4]), .Y(n370) );
  INVX4 U358 ( .A(n137), .Y(n240) );
  XNOR2X2 U359 ( .A(n101), .B(n8), .Y(SUM[24]) );
  CLKINVX2 U360 ( .A(n181), .Y(n180) );
  OAI2BB1X2 U361 ( .A0N(n116), .A1N(n86), .B0(n85), .Y(n83) );
  OR2X2 U362 ( .A(B[15]), .B(A[15]), .Y(n385) );
  NAND2XL U363 ( .A(n385), .B(n160), .Y(n17) );
  XNOR2X1 U364 ( .A(n56), .B(n379), .Y(SUM[29]) );
  INVX3 U365 ( .A(n116), .Y(n115) );
  CLKINVXL U366 ( .A(n142), .Y(n241) );
  INVX1 U367 ( .A(n69), .Y(n71) );
  OAI21X2 U368 ( .A0(n210), .A1(n208), .B0(n209), .Y(n207) );
  NAND2X1 U369 ( .A(n43), .B(n42), .Y(n2) );
  AOI21X2 U370 ( .A0(n370), .A1(n215), .B0(n212), .Y(n210) );
  NAND2X1 U371 ( .A(B[4]), .B(A[4]), .Y(n214) );
  NAND2X1 U372 ( .A(B[7]), .B(A[7]), .Y(n201) );
  NOR2X1 U373 ( .A(n151), .B(n148), .Y(n146) );
  OAI21X1 U374 ( .A0(n164), .A1(n170), .B0(n165), .Y(n163) );
  AOI21X1 U375 ( .A0(n388), .A1(n190), .B0(n185), .Y(n183) );
  NOR2X1 U376 ( .A(n126), .B(n121), .Y(n119) );
  INVX1 U377 ( .A(n192), .Y(n190) );
  NAND2X1 U378 ( .A(B[27]), .B(A[27]), .Y(n75) );
  NOR2X1 U379 ( .A(B[30]), .B(A[30]), .Y(n41) );
  NAND2BXL U380 ( .AN(n224), .B(n225), .Y(n31) );
  OAI21X1 U381 ( .A0(n115), .A1(n393), .B0(n96), .Y(n94) );
  CLKINVXL U382 ( .A(n169), .Y(n246) );
  OAI21X1 U383 ( .A0(n71), .A1(n61), .B0(n64), .Y(n60) );
  NOR2X2 U384 ( .A(B[23]), .B(A[23]), .Y(n110) );
  NAND2X1 U385 ( .A(n242), .B(n149), .Y(n15) );
  AOI21X1 U386 ( .A0(n52), .A1(n69), .B0(n53), .Y(n51) );
  AOI21X1 U387 ( .A0(n48), .A1(n116), .B0(n49), .Y(n47) );
  NAND2X1 U388 ( .A(B[19]), .B(A[19]), .Y(n138) );
  INVX1 U389 ( .A(n187), .Y(n185) );
  INVX2 U390 ( .A(n35), .Y(n378) );
  NAND2X2 U391 ( .A(B[28]), .B(A[28]), .Y(n64) );
  NAND2X1 U392 ( .A(B[30]), .B(A[30]), .Y(n42) );
  OR2X1 U393 ( .A(B[0]), .B(A[0]), .Y(n381) );
  INVX1 U394 ( .A(n160), .Y(n158) );
  CLKINVXL U395 ( .A(n148), .Y(n242) );
  CLKINVXL U396 ( .A(n126), .Y(n239) );
  XOR2X4 U397 ( .A(n139), .B(n372), .Y(SUM[19]) );
  NAND2X4 U398 ( .A(n240), .B(n138), .Y(n372) );
  NAND2XL U399 ( .A(n243), .B(n152), .Y(n16) );
  CLKINVXL U400 ( .A(n143), .Y(n141) );
  NOR2X2 U401 ( .A(B[19]), .B(A[19]), .Y(n137) );
  NAND2X2 U402 ( .A(n394), .B(n131), .Y(n117) );
  OAI2BB1X1 U403 ( .A0N(n116), .A1N(n237), .B0(n114), .Y(n112) );
  XOR2X1 U404 ( .A(n115), .B(n383), .Y(SUM[22]) );
  OAI2BB1X1 U405 ( .A0N(n116), .A1N(n104), .B0(n103), .Y(n101) );
  NAND2XL U406 ( .A(n97), .B(n100), .Y(n8) );
  NAND2XL U407 ( .A(n238), .B(n122), .Y(n373) );
  XOR2X1 U408 ( .A(n177), .B(n374), .Y(SUM[12]) );
  AND2X1 U409 ( .A(n247), .B(n176), .Y(n374) );
  CLKINVXL U410 ( .A(n100), .Y(n98) );
  NAND2XL U411 ( .A(n248), .B(n179), .Y(n21) );
  CLKINVXL U412 ( .A(n178), .Y(n248) );
  CLKINVXL U413 ( .A(n99), .Y(n97) );
  XOR2X1 U414 ( .A(n193), .B(n384), .Y(SUM[9]) );
  XOR2X1 U415 ( .A(n199), .B(n375), .Y(SUM[8]) );
  AND2X1 U416 ( .A(n387), .B(n198), .Y(n375) );
  XNOR2X1 U417 ( .A(n188), .B(n376), .Y(SUM[10]) );
  AND2X1 U418 ( .A(n388), .B(n187), .Y(n376) );
  AOI2BB1X1 U419 ( .A0N(n47), .A1N(n34), .B0(n378), .Y(SUM[32]) );
  NAND2XL U420 ( .A(n68), .B(n52), .Y(n50) );
  CLKINVXL U421 ( .A(n170), .Y(n168) );
  NAND2X2 U422 ( .A(B[22]), .B(A[22]), .Y(n114) );
  NAND2BX1 U423 ( .AN(n74), .B(n75), .Y(n5) );
  NAND2XL U424 ( .A(B[23]), .B(A[23]), .Y(n111) );
  NAND2XL U425 ( .A(B[12]), .B(A[12]), .Y(n176) );
  NAND2XL U426 ( .A(B[8]), .B(A[8]), .Y(n198) );
  NAND2BX1 U427 ( .AN(n216), .B(n217), .Y(n29) );
  XNOR2X4 U428 ( .A(n40), .B(n380), .Y(SUM[31]) );
  NAND2X1 U429 ( .A(n390), .B(n39), .Y(n380) );
  NAND2XL U430 ( .A(n370), .B(n214), .Y(n28) );
  NAND2BX1 U431 ( .AN(n200), .B(n201), .Y(n25) );
  XNOR2XL U432 ( .A(n26), .B(n207), .Y(SUM[6]) );
  NAND2BX1 U433 ( .AN(n208), .B(n209), .Y(n27) );
  OR2X2 U434 ( .A(B[6]), .B(A[6]), .Y(n392) );
  NAND2XL U435 ( .A(B[6]), .B(A[6]), .Y(n206) );
  NAND2XL U436 ( .A(B[2]), .B(A[2]), .Y(n222) );
  NAND2XL U437 ( .A(n391), .B(n222), .Y(n30) );
  INVX2 U438 ( .A(n154), .Y(n153) );
  XNOR2X2 U439 ( .A(n150), .B(n15), .Y(SUM[17]) );
  INVX2 U440 ( .A(n194), .Y(n193) );
  NOR2X1 U441 ( .A(n142), .B(n137), .Y(n131) );
  NOR2X1 U442 ( .A(n133), .B(n126), .Y(n124) );
  XOR2X1 U443 ( .A(n144), .B(n382), .Y(SUM[18]) );
  AND2X1 U444 ( .A(n241), .B(n143), .Y(n382) );
  XOR2X1 U445 ( .A(n161), .B(n17), .Y(SUM[15]) );
  INVX2 U446 ( .A(n172), .Y(n171) );
  CLKINVXL U447 ( .A(n132), .Y(n134) );
  INVX2 U448 ( .A(n164), .Y(n245) );
  XOR2X1 U449 ( .A(n153), .B(n16), .Y(SUM[16]) );
  CLKINVXL U450 ( .A(n151), .Y(n243) );
  NOR2X2 U451 ( .A(B[20]), .B(A[20]), .Y(n126) );
  OAI21X2 U452 ( .A0(n92), .A1(n100), .B0(n93), .Y(n91) );
  NAND2X1 U453 ( .A(n236), .B(n111), .Y(n9) );
  INVX2 U454 ( .A(n110), .Y(n236) );
  CLKINVXL U455 ( .A(n92), .Y(n234) );
  OAI21X1 U456 ( .A0(n110), .A1(n114), .B0(n111), .Y(n105) );
  NAND2X1 U457 ( .A(n237), .B(n114), .Y(n383) );
  NAND2X2 U458 ( .A(B[16]), .B(A[16]), .Y(n152) );
  AOI21X1 U459 ( .A0(n199), .A1(n387), .B0(n196), .Y(n194) );
  INVX2 U460 ( .A(n198), .Y(n196) );
  AND2X1 U461 ( .A(n389), .B(n192), .Y(n384) );
  NAND2XL U462 ( .A(n86), .B(n68), .Y(n66) );
  NAND2X1 U463 ( .A(B[18]), .B(A[18]), .Y(n143) );
  NOR2X1 U464 ( .A(B[14]), .B(A[14]), .Y(n164) );
  NOR2X1 U465 ( .A(B[18]), .B(A[18]), .Y(n142) );
  NAND2X1 U466 ( .A(B[17]), .B(A[17]), .Y(n149) );
  CLKINVXL U467 ( .A(n113), .Y(n237) );
  NAND2X1 U468 ( .A(B[15]), .B(A[15]), .Y(n160) );
  XOR2X1 U469 ( .A(n171), .B(n386), .Y(SUM[13]) );
  AND2X1 U470 ( .A(n246), .B(n170), .Y(n386) );
  NAND2X1 U471 ( .A(n43), .B(n390), .Y(n34) );
  NAND2X1 U472 ( .A(B[14]), .B(A[14]), .Y(n165) );
  OAI21XL U473 ( .A0(n180), .A1(n178), .B0(n179), .Y(n177) );
  INVX2 U474 ( .A(n175), .Y(n247) );
  NOR2X2 U475 ( .A(A[21]), .B(B[21]), .Y(n121) );
  NAND2X1 U476 ( .A(n79), .B(n82), .Y(n6) );
  NAND2X1 U477 ( .A(B[24]), .B(A[24]), .Y(n100) );
  INVX2 U478 ( .A(n82), .Y(n80) );
  NOR2X1 U479 ( .A(B[24]), .B(A[24]), .Y(n99) );
  OAI21X2 U480 ( .A0(n74), .A1(n82), .B0(n75), .Y(n69) );
  NAND2X1 U481 ( .A(n231), .B(n64), .Y(n4) );
  CLKINVXL U482 ( .A(n61), .Y(n231) );
  NOR2X1 U483 ( .A(B[13]), .B(A[13]), .Y(n169) );
  OAI21XL U484 ( .A0(n54), .A1(n64), .B0(n55), .Y(n53) );
  NAND2X1 U485 ( .A(B[13]), .B(A[13]), .Y(n170) );
  OR2X1 U486 ( .A(B[10]), .B(A[10]), .Y(n388) );
  INVX2 U487 ( .A(n206), .Y(n204) );
  INVX2 U488 ( .A(n214), .Y(n212) );
  CLKINVXL U489 ( .A(n81), .Y(n79) );
  OR2X1 U490 ( .A(B[9]), .B(A[9]), .Y(n389) );
  NAND2X1 U491 ( .A(B[10]), .B(A[10]), .Y(n187) );
  NAND2X1 U492 ( .A(B[9]), .B(A[9]), .Y(n192) );
  NAND2X1 U493 ( .A(n392), .B(n206), .Y(n26) );
  INVX2 U494 ( .A(n41), .Y(n43) );
  INVX2 U495 ( .A(n39), .Y(n37) );
  INVX2 U496 ( .A(n42), .Y(n44) );
  OR2X1 U497 ( .A(n261), .B(n260), .Y(n390) );
  NAND2X1 U498 ( .A(n261), .B(n260), .Y(n39) );
  NOR2X1 U499 ( .A(B[3]), .B(A[3]), .Y(n216) );
  INVX2 U500 ( .A(n222), .Y(n220) );
  NAND2X1 U501 ( .A(B[3]), .B(A[3]), .Y(n217) );
  NOR2X1 U502 ( .A(B[5]), .B(A[5]), .Y(n208) );
  NAND2X1 U503 ( .A(B[5]), .B(A[5]), .Y(n209) );
  INVX2 U504 ( .A(A[32]), .Y(n261) );
  INVX2 U505 ( .A(B[32]), .Y(n260) );
  NAND2XL U506 ( .A(B[1]), .B(A[1]), .Y(n225) );
  NAND2X1 U507 ( .A(B[0]), .B(A[0]), .Y(n227) );
  NOR2X1 U508 ( .A(B[22]), .B(A[22]), .Y(n113) );
  NAND2XL U509 ( .A(n104), .B(n97), .Y(n393) );
  OAI21X1 U510 ( .A0(n115), .A1(n66), .B0(n67), .Y(n65) );
  OAI21XL U511 ( .A0(n85), .A1(n50), .B0(n51), .Y(n49) );
  NOR2X4 U512 ( .A(B[28]), .B(A[28]), .Y(n61) );
  NAND2X1 U513 ( .A(n239), .B(n395), .Y(n12) );
  NOR2X1 U514 ( .A(n126), .B(n121), .Y(n394) );
  AOI21X1 U515 ( .A0(n144), .A1(n124), .B0(n125), .Y(n123) );
  CLKINVXL U516 ( .A(n131), .Y(n133) );
  XNOR2X1 U517 ( .A(n28), .B(n215), .Y(SUM[4]) );
  NAND2X1 U518 ( .A(A[21]), .B(B[21]), .Y(n122) );
  NAND2XL U519 ( .A(B[20]), .B(A[20]), .Y(n129) );
  INVX2 U520 ( .A(n105), .Y(n103) );
  NOR2X4 U521 ( .A(n81), .B(n74), .Y(n68) );
  NAND2XL U522 ( .A(n59), .B(n86), .Y(n57) );
  NAND2XL U523 ( .A(B[20]), .B(A[20]), .Y(n395) );
  OAI21X4 U524 ( .A0(n117), .A1(n145), .B0(n118), .Y(n116) );
  OAI21X2 U525 ( .A0(n153), .A1(n151), .B0(n152), .Y(n150) );
  OAI21X1 U526 ( .A0(n224), .A1(n227), .B0(n225), .Y(n223) );
  INVX4 U527 ( .A(n145), .Y(n144) );
  AOI21X4 U528 ( .A0(n154), .A1(n146), .B0(n147), .Y(n145) );
  AOI21X4 U529 ( .A0(n144), .A1(n241), .B0(n141), .Y(n139) );
  OAI21XL U530 ( .A0(n115), .A1(n57), .B0(n58), .Y(n56) );
  OAI21XL U531 ( .A0(n115), .A1(n77), .B0(n78), .Y(n76) );
  NAND2XL U532 ( .A(n86), .B(n79), .Y(n77) );
  AOI21XL U533 ( .A0(n87), .A1(n79), .B0(n80), .Y(n78) );
  OAI21XL U534 ( .A0(n134), .A1(n126), .B0(n395), .Y(n125) );
  OAI21X1 U535 ( .A0(n129), .A1(n121), .B0(n122), .Y(n120) );
  NOR2X4 U536 ( .A(B[29]), .B(A[29]), .Y(n54) );
  AOI21XL U537 ( .A0(n87), .A1(n59), .B0(n60), .Y(n58) );
  NOR2X4 U538 ( .A(B[27]), .B(A[27]), .Y(n74) );
  AOI21XL U539 ( .A0(n87), .A1(n68), .B0(n69), .Y(n67) );
  XOR2X1 U540 ( .A(n25), .B(n202), .Y(SUM[7]) );
  XOR2X1 U541 ( .A(n27), .B(n210), .Y(SUM[5]) );
endmodule


module PE_DW_mult_tc_17 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n6, n9, n12, n16, n18, n22, n24, n30, n34, n36, n40, n42, n46, n48,
         n51, n52, n53, n55, n56, n57, n59, n60, n61, n62, n64, n66, n67, n68,
         n70, n71, n72, n73, n75, n76, n77, n79, n80, n82, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n103, n105, n106, n107, n108, n109, n110, n114, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n140, n141, n142,
         n143, n144, n145, n148, n149, n151, n154, n155, n156, n157, n158,
         n159, n160, n164, n166, n167, n168, n169, n170, n171, n173, n176,
         n177, n181, n182, n183, n184, n185, n186, n187, n188, n191, n192,
         n193, n194, n196, n199, n200, n201, n203, n204, n205, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n219, n220, n221,
         n222, n224, n227, n228, n229, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n244, n245, n246, n247, n248,
         n249, n251, n254, n255, n256, n257, n259, n260, n261, n262, n264,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n281, n283, n284, n286, n288, n289, n290, n292,
         n294, n295, n296, n297, n298, n300, n302, n303, n304, n305, n307,
         n308, n311, n312, n313, n315, n316, n317, n319, n321, n322, n323,
         n324, n325, n326, n327, n329, n334, n336, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n844, n845, n846, n848, n849, n850, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001;

  AOI21X1 U60 ( .A0(n123), .A1(n89), .B0(n90), .Y(n88) );
  AOI21X1 U72 ( .A0(n123), .A1(n98), .B0(n99), .Y(n97) );
  AOI21X1 U76 ( .A0(n114), .A1(n990), .B0(n103), .Y(n101) );
  AOI21X1 U88 ( .A0(n123), .A1(n989), .B0(n114), .Y(n110) );
  AOI21X1 U118 ( .A0(n160), .A1(n135), .B0(n136), .Y(n134) );
  AOI21X1 U132 ( .A0(n160), .A1(n313), .B0(n151), .Y(n145) );
  NOR2X2 U169 ( .A(n370), .B(n363), .Y(n170) );
  NAND2X4 U175 ( .A(n193), .B(n181), .Y(n53) );
  NOR2X2 U211 ( .A(n399), .B(n410), .Y(n204) );
  NOR2X2 U239 ( .A(n227), .B(n232), .Y(n221) );
  NOR2X2 U251 ( .A(n451), .B(n464), .Y(n232) );
  NOR2X2 U270 ( .A(n477), .B(n488), .Y(n245) );
  NOR2X2 U280 ( .A(n489), .B(n498), .Y(n248) );
  NAND2X4 U281 ( .A(n489), .B(n498), .Y(n249) );
  AOI21X1 U286 ( .A0(n327), .A1(n264), .B0(n259), .Y(n257) );
  NOR2X2 U291 ( .A(n499), .B(n508), .Y(n260) );
  NAND2X4 U300 ( .A(n509), .B(n516), .Y(n266) );
  AOI21X1 U320 ( .A0(n985), .A1(n286), .B0(n281), .Y(n279) );
  AOI21X1 U337 ( .A0(n295), .A1(n988), .B0(n292), .Y(n290) );
  ADDFHX4 U381 ( .A(n367), .B(n365), .CI(n372), .CO(n362), .S(n363) );
  ADDFHX4 U385 ( .A(n382), .B(n373), .CI(n380), .CO(n370), .S(n371) );
  ADDFHX4 U389 ( .A(n392), .B(n390), .CI(n381), .CO(n378), .S(n379) );
  ADDFHX4 U399 ( .A(n403), .B(n412), .CI(n401), .CO(n398), .S(n399) );
  ADDFHX4 U411 ( .A(n427), .B(n438), .CI(n425), .CO(n422), .S(n423) );
  ADDFHX4 U418 ( .A(n441), .B(n452), .CI(n439), .CO(n436), .S(n437) );
  ADDFHX4 U426 ( .A(n455), .B(n466), .CI(n453), .CO(n450), .S(n451) );
  ADDFHX4 U439 ( .A(n481), .B(n490), .CI(n479), .CO(n476), .S(n477) );
  ADDFHX4 U445 ( .A(n493), .B(n500), .CI(n491), .CO(n488), .S(n489) );
  ADDFHX4 U450 ( .A(n503), .B(n510), .CI(n501), .CO(n498), .S(n499) );
  ADDFHX4 U455 ( .A(n513), .B(n518), .CI(n511), .CO(n508), .S(n509) );
  OAI22X1 U475 ( .A0(n48), .A1(n868), .B0(n46), .B1(n708), .Y(n556) );
  OAI22X1 U478 ( .A0(n48), .A1(n693), .B0(n692), .B1(n46), .Y(n338) );
  OAI22X1 U479 ( .A0(n48), .A1(n694), .B0(n693), .B1(n46), .Y(n565) );
  OAI22X1 U480 ( .A0(n48), .A1(n695), .B0(n694), .B1(n46), .Y(n566) );
  OAI22X1 U481 ( .A0(n48), .A1(n696), .B0(n695), .B1(n46), .Y(n567) );
  OAI22X1 U483 ( .A0(n48), .A1(n698), .B0(n697), .B1(n46), .Y(n569) );
  OAI22X1 U484 ( .A0(n48), .A1(n699), .B0(n698), .B1(n46), .Y(n570) );
  OAI22X1 U485 ( .A0(n48), .A1(n700), .B0(n699), .B1(n46), .Y(n571) );
  OAI22X1 U487 ( .A0(n48), .A1(n702), .B0(n701), .B1(n46), .Y(n573) );
  OAI22X1 U488 ( .A0(n48), .A1(n703), .B0(n702), .B1(n46), .Y(n574) );
  OAI22X1 U490 ( .A0(n48), .A1(n705), .B0(n704), .B1(n46), .Y(n576) );
  OAI22X1 U491 ( .A0(n48), .A1(n706), .B0(n705), .B1(n46), .Y(n577) );
  OAI22X1 U514 ( .A0(n42), .A1(n710), .B0(n709), .B1(n40), .Y(n344) );
  OAI22X1 U515 ( .A0(n42), .A1(n711), .B0(n710), .B1(n40), .Y(n581) );
  OAI22X1 U516 ( .A0(n42), .A1(n712), .B0(n711), .B1(n40), .Y(n582) );
  OAI22X1 U517 ( .A0(n42), .A1(n713), .B0(n712), .B1(n40), .Y(n583) );
  OAI22X1 U518 ( .A0(n42), .A1(n714), .B0(n713), .B1(n40), .Y(n584) );
  OAI22X1 U519 ( .A0(n42), .A1(n715), .B0(n714), .B1(n40), .Y(n585) );
  OAI22X1 U524 ( .A0(n42), .A1(n720), .B0(n719), .B1(n40), .Y(n590) );
  OAI22X1 U525 ( .A0(n42), .A1(n721), .B0(n720), .B1(n40), .Y(n591) );
  OAI22X1 U526 ( .A0(n42), .A1(n722), .B0(n721), .B1(n40), .Y(n592) );
  OAI22X1 U527 ( .A0(n42), .A1(n723), .B0(n722), .B1(n40), .Y(n593) );
  OAI22X1 U547 ( .A0(n36), .A1(n870), .B0(n961), .B1(n742), .Y(n558) );
  OAI22X1 U593 ( .A0(n30), .A1(n751), .B0(n750), .B1(n993), .Y(n619) );
  OAI22X1 U619 ( .A0(n24), .A1(n872), .B0(n22), .B1(n776), .Y(n560) );
  OAI22X1 U623 ( .A0(n24), .A1(n762), .B0(n761), .B1(n22), .Y(n629) );
  OAI22X1 U625 ( .A0(n24), .A1(n764), .B0(n763), .B1(n22), .Y(n631) );
  OAI22X1 U628 ( .A0(n24), .A1(n767), .B0(n766), .B1(n22), .Y(n634) );
  OAI22X1 U629 ( .A0(n24), .A1(n768), .B0(n767), .B1(n22), .Y(n635) );
  OAI22X1 U630 ( .A0(n24), .A1(n769), .B0(n768), .B1(n22), .Y(n636) );
  OAI22X1 U632 ( .A0(n24), .A1(n771), .B0(n770), .B1(n22), .Y(n638) );
  OAI22X1 U634 ( .A0(n24), .A1(n773), .B0(n772), .B1(n22), .Y(n640) );
  OAI22X1 U635 ( .A0(n24), .A1(n774), .B0(n773), .B1(n22), .Y(n641) );
  OAI22X1 U658 ( .A0(n18), .A1(n778), .B0(n777), .B1(n16), .Y(n408) );
  OAI22X1 U660 ( .A0(n18), .A1(n780), .B0(n779), .B1(n16), .Y(n646) );
  OAI22X1 U664 ( .A0(n18), .A1(n784), .B0(n783), .B1(n16), .Y(n650) );
  OAI22X1 U666 ( .A0(n18), .A1(n786), .B0(n785), .B1(n16), .Y(n652) );
  OAI22X1 U672 ( .A0(n18), .A1(n792), .B0(n791), .B1(n16), .Y(n658) );
  OAI22X1 U699 ( .A0(n12), .A1(n800), .B0(n799), .B1(n9), .Y(n665) );
  OAI22X1 U708 ( .A0(n12), .A1(n809), .B0(n808), .B1(n9), .Y(n674) );
  OAI22X1 U731 ( .A0(n6), .A1(n813), .B0(n812), .B1(n958), .Y(n678) );
  OAI22X1 U732 ( .A0(n6), .A1(n814), .B0(n813), .B1(n958), .Y(n679) );
  OAI22X1 U733 ( .A0(n6), .A1(n815), .B0(n814), .B1(n958), .Y(n680) );
  OAI22X1 U735 ( .A0(n6), .A1(n817), .B0(n816), .B1(n958), .Y(n682) );
  OAI22X1 U738 ( .A0(n6), .A1(n820), .B0(n819), .B1(n958), .Y(n685) );
  OAI22X1 U739 ( .A0(n6), .A1(n821), .B0(n820), .B1(n958), .Y(n686) );
  OAI22X1 U740 ( .A0(n6), .A1(n822), .B0(n821), .B1(n958), .Y(n687) );
  OAI22X1 U742 ( .A0(n6), .A1(n824), .B0(n823), .B1(n958), .Y(n689) );
  OAI22X1 U743 ( .A0(n6), .A1(n825), .B0(n824), .B1(n958), .Y(n690) );
  NAND2X4 U786 ( .A(n46), .B(n844), .Y(n48) );
  XNOR2X4 U788 ( .A(n1000), .B(a[14]), .Y(n46) );
  NAND2X4 U789 ( .A(n40), .B(n845), .Y(n42) );
  XNOR2X4 U791 ( .A(n999), .B(a[12]), .Y(n40) );
  NAND2X4 U792 ( .A(n960), .B(n846), .Y(n36) );
  NAND2X4 U798 ( .A(n22), .B(n848), .Y(n24) );
  XNOR2X4 U800 ( .A(n996), .B(a[6]), .Y(n22) );
  NAND2X4 U801 ( .A(n16), .B(n849), .Y(n18) );
  XNOR2X4 U803 ( .A(n995), .B(a[4]), .Y(n16) );
  NAND2X4 U804 ( .A(n9), .B(n850), .Y(n12) );
  XNOR2X4 U806 ( .A(n994), .B(a[2]), .Y(n9) );
  NOR2X2 U812 ( .A(n211), .B(n216), .Y(n209) );
  NOR2X2 U813 ( .A(n411), .B(n422), .Y(n211) );
  ADDFHX2 U814 ( .A(n456), .B(n443), .CI(n454), .CO(n438), .S(n439) );
  ADDFHX4 U815 ( .A(n462), .B(n449), .CI(n460), .CO(n442), .S(n443) );
  AOI21X1 U816 ( .A0(n234), .A1(n323), .B0(n231), .Y(n229) );
  OAI21XL U817 ( .A0(n242), .A1(n238), .B0(n239), .Y(n237) );
  OAI21X1 U818 ( .A0(n268), .A1(n256), .B0(n257), .Y(n255) );
  INVX3 U819 ( .A(n959), .Y(n962) );
  INVX4 U820 ( .A(n34), .Y(n959) );
  OAI22X1 U821 ( .A0(n36), .A1(n741), .B0(n740), .B1(n962), .Y(n610) );
  XOR2X1 U822 ( .A(n416), .B(n418), .Y(n943) );
  XOR2X1 U823 ( .A(n414), .B(n943), .Y(n401) );
  NAND2X1 U824 ( .A(n416), .B(n414), .Y(n944) );
  NAND2X1 U825 ( .A(n418), .B(n414), .Y(n945) );
  NAND2X1 U826 ( .A(n418), .B(n416), .Y(n946) );
  NAND3X1 U827 ( .A(n945), .B(n946), .C(n944), .Y(n400) );
  ADDFHX2 U828 ( .A(n617), .B(n603), .CI(n432), .CO(n416), .S(n417) );
  ADDFHX1 U829 ( .A(n430), .B(n421), .CI(n419), .CO(n414), .S(n415) );
  ADDFHX2 U830 ( .A(n402), .B(n400), .CI(n391), .CO(n388), .S(n389) );
  OR2X1 U831 ( .A(n30), .B(n756), .Y(n947) );
  OR2X1 U832 ( .A(n755), .B(n993), .Y(n948) );
  NAND2X4 U833 ( .A(n947), .B(n948), .Y(n624) );
  XNOR2X1 U834 ( .A(b[2]), .B(n998), .Y(n756) );
  ADDFHX2 U835 ( .A(n638), .B(n624), .CI(n507), .CO(n502), .S(n503) );
  AND2X1 U836 ( .A(n51), .B(n142), .Y(n949) );
  NOR2X1 U837 ( .A(n949), .B(n143), .Y(n141) );
  AND2X1 U838 ( .A(n51), .B(n155), .Y(n950) );
  NOR2X1 U839 ( .A(n950), .B(n156), .Y(n154) );
  NOR2XL U840 ( .A(n53), .B(n157), .Y(n155) );
  AND2XL U841 ( .A(n51), .B(n168), .Y(n951) );
  NOR2X1 U842 ( .A(n951), .B(n169), .Y(n167) );
  NOR2XL U843 ( .A(n53), .B(n170), .Y(n168) );
  NOR2XL U844 ( .A(n24), .B(n775), .Y(n952) );
  NOR2XL U845 ( .A(n774), .B(n22), .Y(n953) );
  OR2X4 U846 ( .A(n952), .B(n953), .Y(n642) );
  XNOR2XL U847 ( .A(b[0]), .B(n997), .Y(n775) );
  AND2X1 U848 ( .A(n51), .B(n131), .Y(n954) );
  NOR2X1 U849 ( .A(n954), .B(n132), .Y(n130) );
  ADDFHX1 U850 ( .A(n632), .B(n576), .CI(n618), .CO(n430), .S(n431) );
  XNOR2X1 U851 ( .A(b[3]), .B(n1001), .Y(n704) );
  XNOR2X1 U852 ( .A(b[2]), .B(n1001), .Y(n705) );
  ADDFHX1 U853 ( .A(n557), .B(n664), .CI(n636), .CO(n484), .S(n485) );
  INVX1 U854 ( .A(n434), .Y(n955) );
  CLKINVX2 U855 ( .A(n955), .Y(n956) );
  ADDFHX2 U856 ( .A(n415), .B(n424), .CI(n413), .CO(n410), .S(n411) );
  ADDFHX2 U857 ( .A(n442), .B(n429), .CI(n440), .CO(n424), .S(n425) );
  ADDFHX1 U858 ( .A(n560), .B(n642), .CI(n670), .CO(n532), .S(n533) );
  ADDFHX1 U859 ( .A(n643), .B(n686), .CI(n657), .CO(n538), .S(n539) );
  ADDFHX1 U860 ( .A(n559), .B(n626), .CI(n640), .CO(n520), .S(n521) );
  XNOR2X2 U861 ( .A(n192), .B(n981), .Y(product[21]) );
  OAI21X1 U862 ( .A0(n211), .A1(n219), .B0(n212), .Y(n210) );
  ADDFHX1 U863 ( .A(n575), .B(n956), .CI(n660), .CO(n420), .S(n421) );
  ADDFHX1 U864 ( .A(n662), .B(n606), .CI(n620), .CO(n458), .S(n459) );
  ADDFHX1 U865 ( .A(n621), .B(n663), .CI(n649), .CO(n472), .S(n473) );
  OAI21X2 U866 ( .A0(n227), .A1(n233), .B0(n228), .Y(n222) );
  INVXL U867 ( .A(n956), .Y(n435) );
  XNOR2X1 U868 ( .A(b[7]), .B(n999), .Y(n734) );
  XNOR2X1 U869 ( .A(b[7]), .B(n996), .Y(n785) );
  XNOR2X1 U870 ( .A(b[7]), .B(n997), .Y(n768) );
  OAI22XL U871 ( .A0(n30), .A1(n745), .B0(n744), .B1(n993), .Y(n613) );
  OAI22XL U872 ( .A0(n30), .A1(n747), .B0(n746), .B1(n993), .Y(n615) );
  OAI22XL U873 ( .A0(n30), .A1(n744), .B0(n743), .B1(n993), .Y(n368) );
  OAI22XL U874 ( .A0(n30), .A1(n748), .B0(n747), .B1(n993), .Y(n616) );
  OAI22XL U875 ( .A0(n30), .A1(n749), .B0(n748), .B1(n993), .Y(n617) );
  OAI22XL U876 ( .A0(n30), .A1(n746), .B0(n745), .B1(n993), .Y(n614) );
  OAI22XL U877 ( .A0(n30), .A1(n755), .B0(n754), .B1(n993), .Y(n623) );
  OAI22XL U878 ( .A0(n30), .A1(n750), .B0(n749), .B1(n993), .Y(n618) );
  OAI22XL U879 ( .A0(n30), .A1(n752), .B0(n751), .B1(n993), .Y(n620) );
  OAI22XL U880 ( .A0(n30), .A1(n754), .B0(n753), .B1(n993), .Y(n622) );
  OAI22XL U881 ( .A0(n30), .A1(n871), .B0(n993), .B1(n759), .Y(n559) );
  OAI22XL U882 ( .A0(n30), .A1(n757), .B0(n756), .B1(n993), .Y(n625) );
  OAI22XL U883 ( .A0(n30), .A1(n753), .B0(n752), .B1(n993), .Y(n621) );
  OR2X1 U884 ( .A(n633), .B(n591), .Y(n448) );
  OAI22X2 U885 ( .A0(n24), .A1(n766), .B0(n765), .B1(n22), .Y(n633) );
  XOR2X2 U886 ( .A(a[14]), .B(n1001), .Y(n844) );
  INVX3 U887 ( .A(n867), .Y(n957) );
  INVX8 U888 ( .A(n957), .Y(n958) );
  CLKINVXL U889 ( .A(a[0]), .Y(n867) );
  OAI22X1 U890 ( .A0(n48), .A1(n704), .B0(n703), .B1(n46), .Y(n575) );
  XNOR2X1 U891 ( .A(b[13]), .B(n995), .Y(n796) );
  XNOR2X1 U892 ( .A(b[13]), .B(n996), .Y(n779) );
  XNOR2X1 U893 ( .A(b[13]), .B(n997), .Y(n762) );
  ADDFHX1 U894 ( .A(n635), .B(n607), .CI(n486), .CO(n470), .S(n471) );
  XNOR2X1 U895 ( .A(b[8]), .B(n997), .Y(n767) );
  XNOR2X1 U896 ( .A(b[8]), .B(n998), .Y(n750) );
  XNOR2X1 U897 ( .A(b[8]), .B(n996), .Y(n784) );
  ADDFHX1 U898 ( .A(n558), .B(n610), .CI(n666), .CO(n504), .S(n505) );
  XNOR2X2 U899 ( .A(b[14]), .B(n995), .Y(n795) );
  XNOR2X2 U900 ( .A(b[1]), .B(n999), .Y(n740) );
  XNOR2X1 U901 ( .A(b[1]), .B(n1001), .Y(n706) );
  XNOR2X1 U902 ( .A(b[1]), .B(n1000), .Y(n723) );
  XNOR2X1 U903 ( .A(b[15]), .B(n995), .Y(n794) );
  XNOR2X2 U904 ( .A(b[6]), .B(n994), .Y(n820) );
  XNOR2X2 U905 ( .A(b[6]), .B(n999), .Y(n735) );
  XNOR2X1 U906 ( .A(b[6]), .B(n996), .Y(n786) );
  XNOR2X1 U907 ( .A(b[6]), .B(n995), .Y(n803) );
  CLKINVX3 U908 ( .A(n959), .Y(n960) );
  INVX2 U909 ( .A(n959), .Y(n961) );
  NOR2X1 U910 ( .A(n18), .B(n788), .Y(n967) );
  BUFX8 U911 ( .A(a[7]), .Y(n997) );
  OAI22XL U912 ( .A0(n12), .A1(n795), .B0(n794), .B1(n9), .Y(n434) );
  ADDHXL U913 ( .A(n679), .B(n650), .CO(n486), .S(n487) );
  OAI22XL U914 ( .A0(n24), .A1(n761), .B0(n760), .B1(n22), .Y(n386) );
  XOR2X2 U915 ( .A(n997), .B(a[8]), .Y(n992) );
  XNOR2X2 U916 ( .A(n998), .B(a[10]), .Y(n34) );
  BUFX8 U917 ( .A(a[13]), .Y(n1000) );
  BUFX4 U918 ( .A(a[15]), .Y(n1001) );
  INVX2 U919 ( .A(n245), .Y(n325) );
  INVX2 U920 ( .A(n171), .Y(n173) );
  NAND2X2 U921 ( .A(n399), .B(n410), .Y(n205) );
  ADDFX2 U922 ( .A(n360), .B(n353), .CI(n358), .CO(n350), .S(n351) );
  NAND2X1 U923 ( .A(n356), .B(n351), .Y(n149) );
  NOR2X2 U924 ( .A(n188), .B(n183), .Y(n181) );
  XOR2X1 U925 ( .A(n996), .B(a[4]), .Y(n849) );
  ADDFX1 U926 ( .A(n571), .B(n386), .CI(n628), .CO(n376), .S(n377) );
  ADDFX2 U927 ( .A(n585), .B(n599), .CI(n613), .CO(n374), .S(n375) );
  ADDFX2 U928 ( .A(n584), .B(n570), .CI(n369), .CO(n366), .S(n367) );
  CMPR32X1 U929 ( .A(n600), .B(n572), .C(n396), .CO(n382), .S(n383) );
  ADDFX2 U930 ( .A(n361), .B(n359), .CI(n364), .CO(n356), .S(n357) );
  NOR2X1 U931 ( .A(n356), .B(n351), .Y(n148) );
  ADDFX2 U932 ( .A(n582), .B(n568), .CI(n355), .CO(n352), .S(n353) );
  ADDFX2 U933 ( .A(n354), .B(n567), .CI(n596), .CO(n348), .S(n349) );
  NAND2X2 U934 ( .A(n451), .B(n464), .Y(n233) );
  NAND2XL U935 ( .A(n324), .B(n239), .Y(n70) );
  NAND2X1 U936 ( .A(n159), .B(n313), .Y(n144) );
  NAND2X1 U937 ( .A(n122), .B(n98), .Y(n96) );
  OAI21X1 U938 ( .A0(n158), .A1(n124), .B0(n125), .Y(n123) );
  NOR2X1 U939 ( .A(n241), .B(n238), .Y(n236) );
  NOR2BXL U940 ( .AN(n193), .B(n188), .Y(n186) );
  CLKINVX2 U941 ( .A(n182), .Y(n980) );
  OAI21X1 U942 ( .A0(n183), .A1(n191), .B0(n184), .Y(n182) );
  NOR2X1 U943 ( .A(n350), .B(n347), .Y(n137) );
  ADDFX2 U944 ( .A(n659), .B(n688), .CI(n673), .CO(n544), .S(n545) );
  ADDHXL U945 ( .A(n689), .B(n562), .CO(n546), .S(n547) );
  ADDHXL U946 ( .A(n683), .B(n654), .CO(n522), .S(n523) );
  OR2X1 U947 ( .A(n967), .B(n968), .Y(n654) );
  NOR2X1 U948 ( .A(n787), .B(n16), .Y(n968) );
  OAI22X1 U949 ( .A0(n6), .A1(n826), .B0(n825), .B1(n958), .Y(n691) );
  ADDFX2 U950 ( .A(n561), .B(n672), .CI(n543), .CO(n540), .S(n541) );
  NAND2X1 U951 ( .A(n965), .B(n966), .Y(n684) );
  ADDFHX1 U952 ( .A(n639), .B(n653), .CI(n667), .CO(n512), .S(n513) );
  OAI22X1 U953 ( .A0(n24), .A1(n772), .B0(n771), .B1(n22), .Y(n639) );
  ADDFX2 U954 ( .A(n637), .B(n665), .CI(n623), .CO(n494), .S(n495) );
  ADDFHX1 U955 ( .A(n651), .B(n506), .CI(n497), .CO(n492), .S(n493) );
  OAI22X1 U956 ( .A0(n42), .A1(n869), .B0(n40), .B1(n725), .Y(n557) );
  NAND2X1 U957 ( .A(n691), .B(n563), .Y(n307) );
  NOR2X1 U958 ( .A(n690), .B(n675), .Y(n304) );
  OR2X1 U959 ( .A(n531), .B(n536), .Y(n985) );
  ADDFX2 U960 ( .A(n529), .B(n532), .CI(n527), .CO(n524), .S(n525) );
  CMPR32X1 U961 ( .A(n535), .B(n538), .C(n533), .CO(n530), .S(n531) );
  ADDFX2 U962 ( .A(n645), .B(n589), .CI(n631), .CO(n418), .S(n419) );
  ADDFX2 U963 ( .A(n604), .B(n646), .CI(n435), .CO(n432), .S(n433) );
  ADDFX2 U964 ( .A(n634), .B(n463), .CI(n474), .CO(n456), .S(n457) );
  ADDFX2 U965 ( .A(n590), .B(n448), .CI(n446), .CO(n428), .S(n429) );
  XNOR2X1 U966 ( .A(n633), .B(n591), .Y(n449) );
  NOR2X1 U967 ( .A(n525), .B(n530), .Y(n274) );
  ADDFHX1 U968 ( .A(n504), .B(n502), .CI(n495), .CO(n490), .S(n491) );
  ADDFHX1 U969 ( .A(n487), .B(n496), .CI(n494), .CO(n480), .S(n481) );
  ADDFX2 U970 ( .A(n475), .B(n484), .CI(n473), .CO(n468), .S(n469) );
  ADDFX2 U971 ( .A(n482), .B(n471), .CI(n480), .CO(n466), .S(n467) );
  ADDFX2 U972 ( .A(n472), .B(n470), .CI(n459), .CO(n454), .S(n455) );
  ADDFX2 U973 ( .A(n586), .B(n614), .CI(n387), .CO(n384), .S(n385) );
  ADDFX2 U974 ( .A(n629), .B(n587), .CI(n601), .CO(n394), .S(n395) );
  ADDFX2 U975 ( .A(n420), .B(n405), .CI(n407), .CO(n402), .S(n403) );
  ADDFHX1 U976 ( .A(n461), .B(n457), .CI(n468), .CO(n452), .S(n453) );
  ADDFX2 U977 ( .A(n458), .B(n447), .CI(n445), .CO(n440), .S(n441) );
  ADDFX2 U978 ( .A(n428), .B(n417), .CI(n426), .CO(n412), .S(n413) );
  ADDFX2 U979 ( .A(n444), .B(n433), .CI(n431), .CO(n426), .S(n427) );
  INVX2 U980 ( .A(n248), .Y(n326) );
  ADDFHX1 U981 ( .A(n469), .B(n478), .CI(n467), .CO(n464), .S(n465) );
  XNOR2X1 U982 ( .A(n247), .B(n71), .Y(product[13]) );
  OAI21X1 U983 ( .A0(n254), .A1(n248), .B0(n249), .Y(n247) );
  ADDFX2 U984 ( .A(n615), .B(n406), .CI(n404), .CO(n392), .S(n393) );
  ADDFHX1 U985 ( .A(n395), .B(n397), .CI(n393), .CO(n390), .S(n391) );
  ADDFX2 U986 ( .A(n598), .B(n376), .CI(n374), .CO(n364), .S(n365) );
  ADDFX2 U987 ( .A(n384), .B(n377), .CI(n375), .CO(n372), .S(n373) );
  ADDFX2 U988 ( .A(n394), .B(n385), .CI(n383), .CO(n380), .S(n381) );
  ADDFX2 U989 ( .A(n597), .B(n583), .CI(n366), .CO(n358), .S(n359) );
  NAND2X1 U990 ( .A(n327), .B(n984), .Y(n256) );
  NOR2X1 U991 ( .A(n465), .B(n476), .Y(n238) );
  AOI21X1 U992 ( .A0(n325), .A1(n251), .B0(n244), .Y(n242) );
  INVX2 U993 ( .A(n249), .Y(n251) );
  NAND2X1 U994 ( .A(n325), .B(n326), .Y(n241) );
  NAND2X1 U995 ( .A(n322), .B(n228), .Y(n68) );
  NAND2X1 U996 ( .A(n159), .B(n135), .Y(n133) );
  ADDFX2 U997 ( .A(n581), .B(n352), .CI(n349), .CO(n346), .S(n347) );
  XOR2X1 U998 ( .A(n213), .B(n66), .Y(product[18]) );
  XOR2X1 U999 ( .A(n51), .B(n977), .Y(product[19]) );
  XOR2X1 U1000 ( .A(n201), .B(n64), .Y(product[20]) );
  AND2X1 U1001 ( .A(n964), .B(n196), .Y(n192) );
  INVX2 U1002 ( .A(n188), .Y(n317) );
  XOR2X1 U1003 ( .A(n154), .B(n59), .Y(product[25]) );
  NOR2X1 U1004 ( .A(n346), .B(n343), .Y(n128) );
  NOR2X1 U1005 ( .A(n53), .B(n133), .Y(n131) );
  NOR2X1 U1006 ( .A(n53), .B(n120), .Y(n118) );
  XOR2X1 U1007 ( .A(n185), .B(n62), .Y(product[22]) );
  XOR2X1 U1008 ( .A(n176), .B(n61), .Y(product[23]) );
  XNOR2X1 U1009 ( .A(n141), .B(n971), .Y(product[26]) );
  INVX2 U1010 ( .A(n91), .Y(n308) );
  NOR2X1 U1011 ( .A(n53), .B(n87), .Y(n85) );
  AND2X1 U1012 ( .A(n975), .B(n307), .Y(product[1]) );
  OAI22X1 U1013 ( .A0(n18), .A1(n787), .B0(n786), .B1(n16), .Y(n653) );
  ADDFX2 U1014 ( .A(n595), .B(n680), .CI(n609), .CO(n496), .S(n497) );
  OAI22X1 U1015 ( .A0(n12), .A1(n799), .B0(n798), .B1(n9), .Y(n664) );
  INVX2 U1016 ( .A(n979), .Y(n52) );
  OAI2BB1X1 U1017 ( .A0N(n194), .A1N(n181), .B0(n980), .Y(n979) );
  XOR2X1 U1018 ( .A(n229), .B(n68), .Y(product[16]) );
  XOR2X1 U1019 ( .A(n220), .B(n67), .Y(product[17]) );
  INVX2 U1020 ( .A(n235), .Y(n234) );
  AOI21XL U1021 ( .A0(n51), .A1(n177), .B0(n979), .Y(n176) );
  AOI21XL U1022 ( .A0(n51), .A1(n186), .B0(n187), .Y(n185) );
  AOI21X1 U1023 ( .A0(n51), .A1(n319), .B0(n203), .Y(n201) );
  NAND2XL U1024 ( .A(n51), .B(n193), .Y(n964) );
  NOR2X1 U1025 ( .A(n204), .B(n199), .Y(n193) );
  OR2X2 U1026 ( .A(n207), .B(n235), .Y(n969) );
  AOI21X1 U1027 ( .A0(n209), .A1(n222), .B0(n210), .Y(n208) );
  AOI21X1 U1028 ( .A0(n255), .A1(n236), .B0(n237), .Y(n235) );
  OR2X1 U1029 ( .A(n6), .B(n819), .Y(n965) );
  OR2X1 U1030 ( .A(n818), .B(n958), .Y(n966) );
  ADDFHX1 U1031 ( .A(n627), .B(n684), .CI(n641), .CO(n528), .S(n529) );
  INVX3 U1032 ( .A(n266), .Y(n264) );
  XOR2X1 U1033 ( .A(n167), .B(n60), .Y(product[24]) );
  XNOR2X1 U1034 ( .A(b[4]), .B(n996), .Y(n788) );
  XNOR2XL U1035 ( .A(b[5]), .B(n996), .Y(n787) );
  OAI22XL U1036 ( .A0(n6), .A1(n818), .B0(n817), .B1(n958), .Y(n683) );
  NAND2X4 U1037 ( .A(n969), .B(n208), .Y(n51) );
  NAND2XL U1038 ( .A(n209), .B(n221), .Y(n207) );
  NOR2X1 U1039 ( .A(n157), .B(n124), .Y(n122) );
  AOI21X1 U1040 ( .A0(n267), .A1(n984), .B0(n264), .Y(n262) );
  NAND2X1 U1041 ( .A(n315), .B(n983), .Y(n157) );
  INVX2 U1042 ( .A(n148), .Y(n313) );
  INVX1 U1043 ( .A(n288), .Y(n286) );
  OAI21X1 U1044 ( .A0(n304), .A1(n307), .B0(n305), .Y(n303) );
  NAND2XL U1045 ( .A(n547), .B(n674), .Y(n302) );
  XNOR2X1 U1046 ( .A(b[6]), .B(n1001), .Y(n701) );
  INVX2 U1047 ( .A(n170), .Y(n315) );
  AOI21X1 U1048 ( .A0(n214), .A1(n234), .B0(n215), .Y(n213) );
  AOI21X4 U1049 ( .A0(n983), .A1(n173), .B0(n164), .Y(n158) );
  ADDFX1 U1050 ( .A(n521), .B(n526), .CI(n519), .CO(n516), .S(n517) );
  OR2XL U1051 ( .A(n525), .B(n530), .Y(n970) );
  CLKINVX2 U1052 ( .A(n246), .Y(n244) );
  NAND2XL U1053 ( .A(n315), .B(n171), .Y(n61) );
  CLKINVXL U1054 ( .A(n53), .Y(n177) );
  NAND2XL U1055 ( .A(n983), .B(n166), .Y(n60) );
  AOI21X1 U1056 ( .A0(n126), .A1(n151), .B0(n127), .Y(n125) );
  NOR2X1 U1057 ( .A(n137), .B(n128), .Y(n126) );
  NAND2X1 U1058 ( .A(n690), .B(n675), .Y(n305) );
  OR2X1 U1059 ( .A(n691), .B(n563), .Y(n975) );
  ADDFX2 U1060 ( .A(n622), .B(n594), .CI(n608), .CO(n482), .S(n483) );
  CMPR22X1 U1061 ( .A(n677), .B(n648), .CO(n462), .S(n463) );
  NAND2BX1 U1062 ( .AN(b[0]), .B(n1001), .Y(n708) );
  OAI22XL U1063 ( .A0(n6), .A1(n823), .B0(n822), .B1(n958), .Y(n688) );
  ADDFX2 U1064 ( .A(n574), .B(n588), .CI(n616), .CO(n404), .S(n405) );
  ADDFX1 U1065 ( .A(n573), .B(n408), .CI(n644), .CO(n396), .S(n397) );
  XNOR2XL U1066 ( .A(b[6]), .B(n997), .Y(n769) );
  XNOR2XL U1067 ( .A(b[5]), .B(n997), .Y(n770) );
  XNOR2XL U1068 ( .A(b[6]), .B(n1000), .Y(n718) );
  NOR2XL U1069 ( .A(n53), .B(n96), .Y(n94) );
  INVX1 U1070 ( .A(n268), .Y(n267) );
  AND2XL U1071 ( .A(n319), .B(n205), .Y(n977) );
  XNOR2X1 U1072 ( .A(n240), .B(n70), .Y(product[14]) );
  NAND2BX1 U1073 ( .AN(n211), .B(n212), .Y(n66) );
  AOI21XL U1074 ( .A0(n234), .A1(n221), .B0(n222), .Y(n220) );
  NAND2BX1 U1075 ( .AN(n199), .B(n200), .Y(n64) );
  OAI21XL U1076 ( .A0(n52), .A1(n157), .B0(n158), .Y(n156) );
  OAI21XL U1077 ( .A0(n52), .A1(n144), .B0(n145), .Y(n143) );
  XOR2X1 U1078 ( .A(n262), .B(n73), .Y(product[11]) );
  CLKINVXL U1079 ( .A(n277), .Y(n276) );
  XNOR2X1 U1080 ( .A(n273), .B(n75), .Y(product[9]) );
  NAND2XL U1081 ( .A(n329), .B(n272), .Y(n75) );
  CLKINVXL U1082 ( .A(n271), .Y(n329) );
  NAND2XL U1083 ( .A(n411), .B(n422), .Y(n212) );
  NAND2XL U1084 ( .A(n316), .B(n184), .Y(n62) );
  XOR2X1 U1085 ( .A(n276), .B(n76), .Y(product[8]) );
  NAND2XL U1086 ( .A(n313), .B(n149), .Y(n59) );
  NAND2XL U1087 ( .A(n389), .B(n398), .Y(n200) );
  INVX2 U1088 ( .A(n149), .Y(n151) );
  NAND2XL U1089 ( .A(n122), .B(n89), .Y(n87) );
  OR2X4 U1090 ( .A(n509), .B(n516), .Y(n984) );
  NAND2X1 U1091 ( .A(n477), .B(n488), .Y(n246) );
  NAND2XL U1092 ( .A(n525), .B(n530), .Y(n275) );
  NAND2XL U1093 ( .A(n499), .B(n508), .Y(n261) );
  AND2X1 U1094 ( .A(n312), .B(n140), .Y(n971) );
  XOR2X1 U1095 ( .A(n130), .B(n57), .Y(product[27]) );
  XOR2X1 U1096 ( .A(n284), .B(n77), .Y(product[7]) );
  AOI21XL U1097 ( .A0(n289), .A1(n987), .B0(n286), .Y(n284) );
  XOR2X1 U1098 ( .A(n106), .B(n55), .Y(product[29]) );
  XOR2X1 U1099 ( .A(n972), .B(n289), .Y(product[6]) );
  AND2X1 U1100 ( .A(n987), .B(n288), .Y(n972) );
  XOR2X1 U1101 ( .A(n117), .B(n56), .Y(product[28]) );
  XOR2XL U1102 ( .A(n80), .B(n298), .Y(product[4]) );
  NAND2XL U1103 ( .A(n334), .B(n297), .Y(n80) );
  CLKINVXL U1104 ( .A(n296), .Y(n334) );
  XOR2XL U1105 ( .A(n973), .B(n303), .Y(product[3]) );
  AND2X1 U1106 ( .A(n986), .B(n302), .Y(n973) );
  XOR2XL U1107 ( .A(n82), .B(n307), .Y(product[2]) );
  CLKINVXL U1108 ( .A(n304), .Y(n336) );
  XNOR2XL U1109 ( .A(n79), .B(n295), .Y(product[5]) );
  OAI21XL U1110 ( .A0(n52), .A1(n133), .B0(n134), .Y(n132) );
  NAND2XL U1111 ( .A(n362), .B(n357), .Y(n166) );
  XOR2X1 U1112 ( .A(n93), .B(n974), .Y(product[30]) );
  NAND2X1 U1113 ( .A(n308), .B(n92), .Y(n974) );
  NOR2X1 U1114 ( .A(n148), .B(n137), .Y(n135) );
  NAND2XL U1115 ( .A(n531), .B(n536), .Y(n283) );
  ADDFHX2 U1116 ( .A(n485), .B(n483), .CI(n492), .CO(n478), .S(n479) );
  ADDFHX1 U1117 ( .A(n522), .B(n515), .CI(n520), .CO(n510), .S(n511) );
  OR2X2 U1118 ( .A(n541), .B(n544), .Y(n988) );
  NAND2XL U1119 ( .A(n541), .B(n544), .Y(n294) );
  NAND2XL U1120 ( .A(n350), .B(n347), .Y(n140) );
  CMPR32X1 U1121 ( .A(n668), .B(n523), .C(n528), .CO(n518), .S(n519) );
  OAI22XL U1122 ( .A0(n12), .A1(n796), .B0(n795), .B1(n9), .Y(n661) );
  OAI22XL U1123 ( .A0(n30), .A1(n758), .B0(n757), .B1(n993), .Y(n626) );
  OAI22XL U1124 ( .A0(n12), .A1(n798), .B0(n797), .B1(n9), .Y(n663) );
  OAI22XL U1125 ( .A0(n6), .A1(n816), .B0(n815), .B1(n958), .Y(n681) );
  CMPR22X1 U1126 ( .A(n681), .B(n652), .CO(n506), .S(n507) );
  CLKINVXL U1127 ( .A(n995), .Y(n874) );
  OAI22XL U1128 ( .A0(n24), .A1(n765), .B0(n764), .B1(n22), .Y(n632) );
  OAI22XL U1129 ( .A0(n24), .A1(n770), .B0(n769), .B1(n22), .Y(n637) );
  XNOR2XL U1130 ( .A(b[0]), .B(n999), .Y(n741) );
  OAI22XL U1131 ( .A0(n6), .A1(n812), .B0(n811), .B1(n958), .Y(n677) );
  OAI22XL U1132 ( .A0(n24), .A1(n763), .B0(n762), .B1(n22), .Y(n630) );
  OAI22XL U1133 ( .A0(n48), .A1(n701), .B0(n700), .B1(n46), .Y(n572) );
  CLKINVXL U1134 ( .A(n777), .Y(n553) );
  OAI22X1 U1135 ( .A0(n6), .A1(n875), .B0(n827), .B1(n958), .Y(n563) );
  CLKINVXL U1136 ( .A(n994), .Y(n875) );
  NAND2BXL U1137 ( .AN(b[0]), .B(n994), .Y(n827) );
  CLKINVXL U1138 ( .A(n794), .Y(n554) );
  NAND2BXL U1139 ( .AN(b[0]), .B(n997), .Y(n776) );
  OAI22XL U1140 ( .A0(n42), .A1(n719), .B0(n718), .B1(n40), .Y(n589) );
  NAND2BXL U1141 ( .AN(b[0]), .B(n1000), .Y(n725) );
  OAI22XL U1142 ( .A0(n42), .A1(n718), .B0(n717), .B1(n40), .Y(n588) );
  XNOR2XL U1143 ( .A(b[0]), .B(n995), .Y(n809) );
  NAND2BXL U1144 ( .AN(b[0]), .B(n995), .Y(n810) );
  NAND2BXL U1145 ( .AN(b[0]), .B(n996), .Y(n793) );
  OAI22XL U1146 ( .A0(n42), .A1(n717), .B0(n716), .B1(n40), .Y(n587) );
  INVX1 U1147 ( .A(n386), .Y(n387) );
  OAI22XL U1148 ( .A0(n42), .A1(n716), .B0(n715), .B1(n40), .Y(n586) );
  CLKINVXL U1149 ( .A(n760), .Y(n552) );
  CLKINVXL U1150 ( .A(n998), .Y(n871) );
  CLKINVXL U1151 ( .A(n1000), .Y(n869) );
  CLKINVXL U1152 ( .A(n999), .Y(n870) );
  CLKINVXL U1153 ( .A(n996), .Y(n873) );
  CLKINVXL U1154 ( .A(n1001), .Y(n868) );
  OAI22XL U1155 ( .A0(n48), .A1(n697), .B0(n696), .B1(n46), .Y(n568) );
  NAND2X4 U1156 ( .A(n976), .B(n958), .Y(n6) );
  XOR2X2 U1157 ( .A(n994), .B(a[0]), .Y(n976) );
  XNOR2XL U1158 ( .A(b[15]), .B(n994), .Y(n811) );
  XNOR2X1 U1159 ( .A(b[5]), .B(n1001), .Y(n702) );
  XNOR2X1 U1160 ( .A(b[8]), .B(n1001), .Y(n699) );
  XNOR2XL U1161 ( .A(b[15]), .B(n999), .Y(n726) );
  XNOR2XL U1162 ( .A(b[15]), .B(n1001), .Y(n692) );
  INVX2 U1163 ( .A(n122), .Y(n120) );
  CLKINVXL U1164 ( .A(n227), .Y(n322) );
  OAI21X1 U1165 ( .A0(n199), .A1(n205), .B0(n200), .Y(n194) );
  INVX2 U1166 ( .A(n255), .Y(n254) );
  XOR2X1 U1167 ( .A(n234), .B(n978), .Y(product[15]) );
  AND2X1 U1168 ( .A(n323), .B(n233), .Y(n978) );
  NAND2XL U1169 ( .A(n321), .B(n219), .Y(n67) );
  CLKINVXL U1170 ( .A(n216), .Y(n321) );
  INVX2 U1171 ( .A(n158), .Y(n160) );
  INVX2 U1172 ( .A(n157), .Y(n159) );
  NOR2BXL U1173 ( .AN(n221), .B(n216), .Y(n214) );
  OAI21XL U1174 ( .A0(n224), .A1(n216), .B0(n219), .Y(n215) );
  CLKINVXL U1175 ( .A(n222), .Y(n224) );
  CLKINVXL U1176 ( .A(n232), .Y(n323) );
  OAI21XL U1177 ( .A0(n254), .A1(n241), .B0(n242), .Y(n240) );
  CLKINVXL U1178 ( .A(n238), .Y(n324) );
  CLKINVXL U1179 ( .A(n204), .Y(n319) );
  CLKINVXL U1180 ( .A(n233), .Y(n231) );
  CLKINVXL U1181 ( .A(n205), .Y(n203) );
  OAI21XL U1182 ( .A0(n52), .A1(n96), .B0(n97), .Y(n95) );
  INVX2 U1183 ( .A(n101), .Y(n99) );
  OAI21XL U1184 ( .A0(n52), .A1(n87), .B0(n88), .Y(n86) );
  INVX2 U1185 ( .A(n261), .Y(n259) );
  AOI21X1 U1186 ( .A0(n269), .A1(n277), .B0(n270), .Y(n268) );
  OAI21X1 U1187 ( .A0(n271), .A1(n275), .B0(n272), .Y(n270) );
  NOR2X1 U1188 ( .A(n271), .B(n274), .Y(n269) );
  NAND2X1 U1189 ( .A(n313), .B(n126), .Y(n124) );
  INVX2 U1190 ( .A(n166), .Y(n164) );
  CLKINVXL U1191 ( .A(n183), .Y(n316) );
  NAND2XL U1192 ( .A(n327), .B(n261), .Y(n73) );
  AND2X1 U1193 ( .A(n317), .B(n191), .Y(n981) );
  NAND2XL U1194 ( .A(n325), .B(n246), .Y(n71) );
  NAND2X2 U1195 ( .A(n437), .B(n450), .Y(n228) );
  OAI21XL U1196 ( .A0(n52), .A1(n170), .B0(n171), .Y(n169) );
  OAI21X1 U1197 ( .A0(n276), .A1(n274), .B0(n275), .Y(n273) );
  NAND2X1 U1198 ( .A(n970), .B(n275), .Y(n76) );
  XOR2X1 U1199 ( .A(n254), .B(n72), .Y(product[12]) );
  NAND2XL U1200 ( .A(n326), .B(n249), .Y(n72) );
  OAI21XL U1201 ( .A0(n52), .A1(n120), .B0(n121), .Y(n119) );
  CLKINVXL U1202 ( .A(n123), .Y(n121) );
  XOR2X1 U1203 ( .A(n267), .B(n982), .Y(product[10]) );
  AND2X1 U1204 ( .A(n984), .B(n266), .Y(n982) );
  NAND2X1 U1205 ( .A(n465), .B(n476), .Y(n239) );
  OAI21XL U1206 ( .A0(n196), .A1(n188), .B0(n191), .Y(n187) );
  CLKINVXL U1207 ( .A(n194), .Y(n196) );
  INVX2 U1208 ( .A(n100), .Y(n98) );
  OAI21XL U1209 ( .A0(n140), .A1(n128), .B0(n129), .Y(n127) );
  OAI21X1 U1210 ( .A0(n101), .A1(n91), .B0(n92), .Y(n90) );
  OAI21X1 U1211 ( .A0(n278), .A1(n290), .B0(n279), .Y(n277) );
  NAND2X1 U1212 ( .A(n985), .B(n987), .Y(n278) );
  INVX2 U1213 ( .A(n283), .Y(n281) );
  OAI21XL U1214 ( .A0(n52), .A1(n109), .B0(n110), .Y(n108) );
  NAND2X1 U1215 ( .A(n990), .B(n105), .Y(n55) );
  NOR2XL U1216 ( .A(n53), .B(n109), .Y(n107) );
  OR2X4 U1217 ( .A(n362), .B(n357), .Y(n983) );
  NAND2X1 U1218 ( .A(n311), .B(n129), .Y(n57) );
  CLKINVXL U1219 ( .A(n128), .Y(n311) );
  OAI21XL U1220 ( .A0(n149), .A1(n137), .B0(n140), .Y(n136) );
  CLKINVXL U1221 ( .A(n137), .Y(n312) );
  INVX2 U1222 ( .A(n294), .Y(n292) );
  AOI21X1 U1223 ( .A0(n986), .A1(n303), .B0(n300), .Y(n298) );
  INVX2 U1224 ( .A(n302), .Y(n300) );
  OAI21X1 U1225 ( .A0(n298), .A1(n296), .B0(n297), .Y(n295) );
  NAND2X2 U1226 ( .A(n370), .B(n363), .Y(n171) );
  NAND2X1 U1227 ( .A(n122), .B(n989), .Y(n109) );
  NOR2X1 U1228 ( .A(n517), .B(n524), .Y(n271) );
  NAND2X1 U1229 ( .A(n989), .B(n116), .Y(n56) );
  NAND2X2 U1230 ( .A(n379), .B(n388), .Y(n191) );
  NAND2X1 U1231 ( .A(n985), .B(n283), .Y(n77) );
  NAND2X1 U1232 ( .A(n378), .B(n371), .Y(n184) );
  NAND2X1 U1233 ( .A(n517), .B(n524), .Y(n272) );
  NAND2X1 U1234 ( .A(n336), .B(n305), .Y(n82) );
  NAND2X1 U1235 ( .A(n988), .B(n294), .Y(n79) );
  INVX2 U1236 ( .A(n105), .Y(n103) );
  INVX2 U1237 ( .A(n116), .Y(n114) );
  NAND2X1 U1238 ( .A(n989), .B(n990), .Y(n100) );
  NOR2X1 U1239 ( .A(n100), .B(n91), .Y(n89) );
  ADDFHX1 U1240 ( .A(n514), .B(n512), .CI(n505), .CO(n500), .S(n501) );
  OR2X2 U1241 ( .A(n547), .B(n674), .Y(n986) );
  NOR2X1 U1242 ( .A(n545), .B(n546), .Y(n296) );
  NAND2X1 U1243 ( .A(n537), .B(n540), .Y(n288) );
  OR2X1 U1244 ( .A(n537), .B(n540), .Y(n987) );
  NAND2XL U1245 ( .A(n346), .B(n343), .Y(n129) );
  NAND2X1 U1246 ( .A(n545), .B(n546), .Y(n297) );
  NAND2X1 U1247 ( .A(n342), .B(n341), .Y(n116) );
  OR2X1 U1248 ( .A(n342), .B(n341), .Y(n989) );
  OR2X1 U1249 ( .A(n340), .B(n339), .Y(n990) );
  INVX2 U1250 ( .A(n338), .Y(n339) );
  NAND2X1 U1251 ( .A(n340), .B(n339), .Y(n105) );
  NOR2X1 U1252 ( .A(n564), .B(n338), .Y(n91) );
  NAND2X1 U1253 ( .A(n564), .B(n338), .Y(n92) );
  INVX2 U1254 ( .A(n726), .Y(n550) );
  NOR2BXL U1255 ( .AN(b[0]), .B(n40), .Y(n595) );
  ADDFHX1 U1256 ( .A(n647), .B(n577), .CI(n605), .CO(n444), .S(n445) );
  ADDFX1 U1257 ( .A(n669), .B(n655), .CI(n534), .CO(n526), .S(n527) );
  ADDFHX1 U1258 ( .A(n556), .B(n578), .CI(n592), .CO(n460), .S(n461) );
  OAI22XL U1259 ( .A0(n48), .A1(n707), .B0(n706), .B1(n46), .Y(n578) );
  ADDFX2 U1260 ( .A(n579), .B(n678), .CI(n593), .CO(n474), .S(n475) );
  NOR2BXL U1261 ( .AN(b[0]), .B(n46), .Y(n579) );
  OAI2BB1X1 U1262 ( .A0N(n958), .A1N(n6), .B0(n555), .Y(n676) );
  ADDFHX1 U1263 ( .A(n611), .B(n682), .CI(n625), .CO(n514), .S(n515) );
  ADDFHX1 U1264 ( .A(n602), .B(n630), .CI(n409), .CO(n406), .S(n407) );
  INVX1 U1265 ( .A(n368), .Y(n369) );
  OAI2BB1X1 U1266 ( .A0N(n22), .A1N(n24), .B0(n552), .Y(n628) );
  ADDFX2 U1267 ( .A(n566), .B(n345), .CI(n348), .CO(n342), .S(n343) );
  INVX1 U1268 ( .A(n344), .Y(n345) );
  NAND2BXL U1269 ( .AN(b[0]), .B(n999), .Y(n742) );
  INVX2 U1270 ( .A(n992), .Y(n993) );
  CLKINVXL U1271 ( .A(n354), .Y(n355) );
  OAI22XL U1272 ( .A0(n42), .A1(n724), .B0(n723), .B1(n40), .Y(n594) );
  ADDFX1 U1273 ( .A(n569), .B(n368), .CI(n612), .CO(n360), .S(n361) );
  OAI2BB1X1 U1274 ( .A0N(n993), .A1N(n30), .B0(n551), .Y(n612) );
  INVX2 U1275 ( .A(n743), .Y(n551) );
  NAND2BX1 U1276 ( .AN(b[0]), .B(n998), .Y(n759) );
  ADDHXL U1277 ( .A(n685), .B(n656), .CO(n534), .S(n535) );
  NOR2BXL U1278 ( .AN(b[0]), .B(n993), .Y(n627) );
  ADDFX2 U1279 ( .A(n671), .B(n542), .CI(n539), .CO(n536), .S(n537) );
  NOR2BXL U1280 ( .AN(b[0]), .B(n22), .Y(n643) );
  XNOR2X1 U1281 ( .A(b[0]), .B(n998), .Y(n758) );
  ADDHXL U1282 ( .A(n687), .B(n658), .CO(n542), .S(n543) );
  ADDFX2 U1283 ( .A(n344), .B(n565), .CI(n580), .CO(n340), .S(n341) );
  OAI2BB1X1 U1284 ( .A0N(n40), .A1N(n42), .B0(n549), .Y(n580) );
  INVX2 U1285 ( .A(n709), .Y(n549) );
  NOR2BXL U1286 ( .AN(b[0]), .B(n9), .Y(n675) );
  INVX2 U1287 ( .A(n811), .Y(n555) );
  INVX2 U1288 ( .A(n997), .Y(n872) );
  NOR2BXL U1289 ( .AN(b[0]), .B(n958), .Y(product[0]) );
  OAI2BB1X1 U1290 ( .A0N(n46), .A1N(n48), .B0(n548), .Y(n564) );
  INVX2 U1291 ( .A(n692), .Y(n548) );
  XOR2X1 U1292 ( .A(n999), .B(a[10]), .Y(n846) );
  BUFX12 U1293 ( .A(a[9]), .Y(n998) );
  XOR2X1 U1294 ( .A(n997), .B(a[6]), .Y(n848) );
  BUFX12 U1295 ( .A(a[5]), .Y(n996) );
  XOR2X1 U1296 ( .A(n995), .B(a[2]), .Y(n850) );
  BUFX12 U1297 ( .A(a[1]), .Y(n994) );
  BUFX12 U1298 ( .A(a[3]), .Y(n995) );
  XOR2X1 U1299 ( .A(n1000), .B(a[12]), .Y(n845) );
  BUFX12 U1300 ( .A(a[11]), .Y(n999) );
  OR2X4 U1301 ( .A(n992), .B(n991), .Y(n30) );
  XNOR2X1 U1302 ( .A(n998), .B(a[8]), .Y(n991) );
  XNOR2XL U1303 ( .A(b[12]), .B(n994), .Y(n814) );
  XNOR2XL U1304 ( .A(b[10]), .B(n994), .Y(n816) );
  XNOR2XL U1305 ( .A(b[14]), .B(n999), .Y(n727) );
  XNOR2XL U1306 ( .A(b[11]), .B(n994), .Y(n815) );
  XNOR2XL U1307 ( .A(b[14]), .B(n994), .Y(n812) );
  XNOR2XL U1308 ( .A(b[9]), .B(n994), .Y(n817) );
  XNOR2XL U1309 ( .A(b[13]), .B(n994), .Y(n813) );
  XNOR2XL U1310 ( .A(b[15]), .B(n998), .Y(n743) );
  XNOR2XL U1311 ( .A(b[4]), .B(n994), .Y(n822) );
  XNOR2XL U1312 ( .A(b[8]), .B(n994), .Y(n818) );
  XNOR2XL U1313 ( .A(b[4]), .B(n999), .Y(n737) );
  XNOR2XL U1314 ( .A(b[5]), .B(n999), .Y(n736) );
  XNOR2XL U1315 ( .A(b[3]), .B(n994), .Y(n823) );
  XNOR2XL U1316 ( .A(b[12]), .B(n996), .Y(n780) );
  XNOR2XL U1317 ( .A(b[12]), .B(n999), .Y(n729) );
  XNOR2XL U1318 ( .A(b[12]), .B(n995), .Y(n797) );
  XNOR2XL U1319 ( .A(b[14]), .B(n998), .Y(n744) );
  XNOR2XL U1320 ( .A(b[3]), .B(n996), .Y(n789) );
  XNOR2XL U1321 ( .A(b[5]), .B(n994), .Y(n821) );
  XNOR2XL U1322 ( .A(b[6]), .B(n998), .Y(n752) );
  XNOR2XL U1323 ( .A(b[7]), .B(n994), .Y(n819) );
  XNOR2XL U1324 ( .A(b[10]), .B(n995), .Y(n799) );
  XNOR2XL U1325 ( .A(b[3]), .B(n999), .Y(n738) );
  XNOR2XL U1326 ( .A(b[2]), .B(n999), .Y(n739) );
  XNOR2XL U1327 ( .A(b[11]), .B(n996), .Y(n781) );
  XNOR2XL U1328 ( .A(b[9]), .B(n999), .Y(n732) );
  XNOR2XL U1329 ( .A(b[11]), .B(n995), .Y(n798) );
  XNOR2XL U1330 ( .A(b[11]), .B(n999), .Y(n730) );
  XNOR2XL U1331 ( .A(b[15]), .B(n997), .Y(n760) );
  XNOR2XL U1332 ( .A(b[1]), .B(n998), .Y(n757) );
  XNOR2XL U1333 ( .A(b[5]), .B(n998), .Y(n753) );
  XNOR2XL U1334 ( .A(b[4]), .B(n997), .Y(n771) );
  XNOR2XL U1335 ( .A(b[7]), .B(n998), .Y(n751) );
  XNOR2XL U1336 ( .A(b[9]), .B(n995), .Y(n800) );
  XNOR2XL U1337 ( .A(b[8]), .B(n999), .Y(n733) );
  XNOR2XL U1338 ( .A(b[2]), .B(n994), .Y(n824) );
  XNOR2XL U1339 ( .A(b[1]), .B(n997), .Y(n774) );
  XNOR2XL U1340 ( .A(b[4]), .B(n1000), .Y(n720) );
  XNOR2XL U1341 ( .A(b[11]), .B(n997), .Y(n764) );
  XNOR2XL U1342 ( .A(b[3]), .B(n998), .Y(n755) );
  XNOR2XL U1343 ( .A(b[2]), .B(n1000), .Y(n722) );
  XNOR2XL U1344 ( .A(b[10]), .B(n997), .Y(n765) );
  XNOR2XL U1345 ( .A(b[3]), .B(n997), .Y(n772) );
  XNOR2XL U1346 ( .A(b[3]), .B(n1000), .Y(n721) );
  XNOR2XL U1347 ( .A(b[10]), .B(n996), .Y(n782) );
  XNOR2XL U1348 ( .A(b[15]), .B(n996), .Y(n777) );
  XNOR2XL U1349 ( .A(b[4]), .B(n1001), .Y(n703) );
  XNOR2XL U1350 ( .A(b[14]), .B(n997), .Y(n761) );
  XNOR2XL U1351 ( .A(b[12]), .B(n997), .Y(n763) );
  XNOR2XL U1352 ( .A(b[9]), .B(n996), .Y(n783) );
  XNOR2XL U1353 ( .A(b[13]), .B(n998), .Y(n745) );
  XNOR2XL U1354 ( .A(b[4]), .B(n998), .Y(n754) );
  XNOR2XL U1355 ( .A(b[9]), .B(n997), .Y(n766) );
  XNOR2XL U1356 ( .A(b[7]), .B(n1000), .Y(n717) );
  XNOR2XL U1357 ( .A(b[2]), .B(n996), .Y(n790) );
  XNOR2XL U1358 ( .A(b[5]), .B(n995), .Y(n804) );
  XNOR2XL U1359 ( .A(b[9]), .B(n1000), .Y(n715) );
  XNOR2XL U1360 ( .A(b[1]), .B(n994), .Y(n825) );
  XNOR2XL U1361 ( .A(b[8]), .B(n995), .Y(n801) );
  XNOR2XL U1362 ( .A(b[14]), .B(n996), .Y(n778) );
  XNOR2XL U1363 ( .A(b[12]), .B(n998), .Y(n746) );
  XNOR2XL U1364 ( .A(b[9]), .B(n1001), .Y(n698) );
  XNOR2XL U1365 ( .A(b[2]), .B(n995), .Y(n807) );
  XNOR2XL U1366 ( .A(b[1]), .B(n996), .Y(n791) );
  XNOR2XL U1367 ( .A(b[8]), .B(n1000), .Y(n716) );
  XNOR2XL U1368 ( .A(b[11]), .B(n1000), .Y(n713) );
  XNOR2XL U1369 ( .A(b[4]), .B(n995), .Y(n805) );
  XNOR2XL U1370 ( .A(b[7]), .B(n1001), .Y(n700) );
  XNOR2XL U1371 ( .A(b[10]), .B(n1000), .Y(n714) );
  XNOR2XL U1372 ( .A(b[2]), .B(n997), .Y(n773) );
  XNOR2XL U1373 ( .A(b[5]), .B(n1000), .Y(n719) );
  XNOR2XL U1374 ( .A(b[11]), .B(n1001), .Y(n696) );
  XNOR2XL U1375 ( .A(b[1]), .B(n995), .Y(n808) );
  XNOR2XL U1376 ( .A(b[12]), .B(n1001), .Y(n695) );
  XNOR2XL U1377 ( .A(b[7]), .B(n995), .Y(n802) );
  XNOR2XL U1378 ( .A(b[10]), .B(n1001), .Y(n697) );
  XNOR2XL U1379 ( .A(b[3]), .B(n995), .Y(n806) );
  XNOR2XL U1380 ( .A(b[13]), .B(n1000), .Y(n711) );
  XNOR2XL U1381 ( .A(b[12]), .B(n1000), .Y(n712) );
  XNOR2XL U1382 ( .A(b[10]), .B(n999), .Y(n731) );
  XNOR2XL U1383 ( .A(b[10]), .B(n998), .Y(n748) );
  XNOR2XL U1384 ( .A(b[9]), .B(n998), .Y(n749) );
  XNOR2XL U1385 ( .A(b[13]), .B(n999), .Y(n728) );
  XNOR2XL U1386 ( .A(b[11]), .B(n998), .Y(n747) );
  XNOR2XL U1387 ( .A(b[15]), .B(n1000), .Y(n709) );
  XNOR2XL U1388 ( .A(b[14]), .B(n1000), .Y(n710) );
  XNOR2XL U1389 ( .A(b[13]), .B(n1001), .Y(n694) );
  XNOR2XL U1390 ( .A(b[14]), .B(n1001), .Y(n693) );
  XNOR2XL U1391 ( .A(b[0]), .B(n1000), .Y(n724) );
  INVX1 U1392 ( .A(n408), .Y(n409) );
  AOI21XL U1393 ( .A0(n51), .A1(n85), .B0(n86), .Y(product[31]) );
  AOI21XL U1394 ( .A0(n51), .A1(n94), .B0(n95), .Y(n93) );
  AOI21XL U1395 ( .A0(n51), .A1(n107), .B0(n108), .Y(n106) );
  AOI21XL U1396 ( .A0(n51), .A1(n118), .B0(n119), .Y(n117) );
  OAI2BB1X1 U1397 ( .A0N(n962), .A1N(n36), .B0(n550), .Y(n596) );
  OAI22XL U1398 ( .A0(n36), .A1(n729), .B0(n728), .B1(n961), .Y(n598) );
  OAI22XL U1399 ( .A0(n36), .A1(n728), .B0(n727), .B1(n961), .Y(n597) );
  OAI22XL U1400 ( .A0(n36), .A1(n731), .B0(n730), .B1(n962), .Y(n600) );
  OAI22XL U1401 ( .A0(n36), .A1(n732), .B0(n731), .B1(n961), .Y(n601) );
  OAI22XL U1402 ( .A0(n36), .A1(n727), .B0(n726), .B1(n962), .Y(n354) );
  OAI22XL U1403 ( .A0(n36), .A1(n730), .B0(n729), .B1(n962), .Y(n599) );
  OAI22XL U1404 ( .A0(n36), .A1(n736), .B0(n735), .B1(n961), .Y(n605) );
  OAI22XL U1405 ( .A0(n36), .A1(n734), .B0(n733), .B1(n961), .Y(n603) );
  OAI22XL U1406 ( .A0(n36), .A1(n739), .B0(n738), .B1(n962), .Y(n608) );
  NOR2BXL U1407 ( .AN(b[0]), .B(n962), .Y(n611) );
  OAI22XL U1408 ( .A0(n36), .A1(n733), .B0(n732), .B1(n961), .Y(n602) );
  OAI22XL U1409 ( .A0(n36), .A1(n740), .B0(n739), .B1(n962), .Y(n609) );
  OAI22XL U1410 ( .A0(n36), .A1(n735), .B0(n734), .B1(n962), .Y(n604) );
  OAI22XL U1411 ( .A0(n36), .A1(n738), .B0(n737), .B1(n961), .Y(n607) );
  OAI22XL U1412 ( .A0(n36), .A1(n737), .B0(n736), .B1(n961), .Y(n606) );
  NOR2X4 U1413 ( .A(n378), .B(n371), .Y(n183) );
  OAI22XL U1414 ( .A0(n12), .A1(n807), .B0(n806), .B1(n9), .Y(n672) );
  OAI22XL U1415 ( .A0(n12), .A1(n808), .B0(n807), .B1(n9), .Y(n673) );
  OAI22XL U1416 ( .A0(n12), .A1(n804), .B0(n803), .B1(n9), .Y(n669) );
  OAI22XL U1417 ( .A0(n12), .A1(n803), .B0(n802), .B1(n9), .Y(n668) );
  OAI2BB1X1 U1418 ( .A0N(n9), .A1N(n12), .B0(n554), .Y(n660) );
  OAI22XL U1419 ( .A0(n12), .A1(n806), .B0(n805), .B1(n9), .Y(n671) );
  OAI22XL U1420 ( .A0(n12), .A1(n802), .B0(n801), .B1(n9), .Y(n667) );
  OAI22XL U1421 ( .A0(n12), .A1(n805), .B0(n804), .B1(n9), .Y(n670) );
  OAI22XL U1422 ( .A0(n12), .A1(n801), .B0(n800), .B1(n9), .Y(n666) );
  OAI22XL U1423 ( .A0(n12), .A1(n874), .B0(n9), .B1(n810), .Y(n562) );
  OAI22XL U1424 ( .A0(n12), .A1(n797), .B0(n796), .B1(n9), .Y(n662) );
  NOR2X4 U1425 ( .A(n389), .B(n398), .Y(n199) );
  NAND2X2 U1426 ( .A(n423), .B(n436), .Y(n219) );
  OAI22X1 U1427 ( .A0(n18), .A1(n782), .B0(n781), .B1(n16), .Y(n648) );
  ADDFHX1 U1428 ( .A(n619), .B(n661), .CI(n676), .CO(n446), .S(n447) );
  OAI2BB1X1 U1429 ( .A0N(n16), .A1N(n18), .B0(n553), .Y(n644) );
  OAI22XL U1430 ( .A0(n18), .A1(n783), .B0(n782), .B1(n16), .Y(n649) );
  OAI22XL U1431 ( .A0(n18), .A1(n779), .B0(n778), .B1(n16), .Y(n645) );
  OAI22XL U1432 ( .A0(n18), .A1(n791), .B0(n790), .B1(n16), .Y(n657) );
  OAI22XL U1433 ( .A0(n18), .A1(n789), .B0(n788), .B1(n16), .Y(n655) );
  NOR2BXL U1434 ( .AN(b[0]), .B(n16), .Y(n659) );
  OAI22XL U1435 ( .A0(n18), .A1(n785), .B0(n784), .B1(n16), .Y(n651) );
  OAI22XL U1436 ( .A0(n18), .A1(n873), .B0(n16), .B1(n793), .Y(n561) );
  OAI22XL U1437 ( .A0(n18), .A1(n790), .B0(n789), .B1(n16), .Y(n656) );
  OAI22XL U1438 ( .A0(n18), .A1(n781), .B0(n780), .B1(n16), .Y(n647) );
  XNOR2XL U1439 ( .A(b[0]), .B(n1001), .Y(n707) );
  NOR2X4 U1440 ( .A(n437), .B(n450), .Y(n227) );
  INVX3 U1441 ( .A(n260), .Y(n327) );
  INVX2 U1442 ( .A(n290), .Y(n289) );
  NOR2XL U1443 ( .A(n53), .B(n144), .Y(n142) );
  NOR2X4 U1444 ( .A(n423), .B(n436), .Y(n216) );
  NOR2X4 U1445 ( .A(n379), .B(n388), .Y(n188) );
  XNOR2X1 U1446 ( .A(b[0]), .B(n996), .Y(n792) );
  XNOR2X1 U1447 ( .A(b[0]), .B(n994), .Y(n826) );
endmodule


module PE_DW_mult_tc_22 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n6, n9, n12, n16, n18, n22, n24, n28, n30, n34, n36, n40, n42, n46,
         n48, n51, n52, n53, n56, n59, n60, n62, n63, n64, n66, n67, n68, n70,
         n71, n72, n73, n75, n76, n77, n79, n80, n81, n82, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n103, n105, n106, n107, n108, n109, n110, n114, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n140, n141, n142,
         n143, n144, n145, n148, n149, n151, n154, n155, n156, n157, n158,
         n159, n160, n164, n166, n167, n168, n169, n170, n171, n176, n177,
         n178, n181, n182, n183, n184, n185, n186, n187, n188, n191, n192,
         n193, n194, n196, n199, n200, n201, n203, n204, n205, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n219, n220, n221,
         n222, n224, n227, n228, n229, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n244, n246, n247, n248, n249,
         n251, n254, n255, n256, n257, n259, n261, n262, n264, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n279,
         n281, n283, n284, n286, n288, n290, n292, n294, n295, n296, n297,
         n298, n300, n302, n303, n304, n305, n307, n308, n311, n312, n313,
         n315, n316, n319, n320, n321, n323, n324, n326, n329, n330, n334,
         n336, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n844, n845, n846, n847,
         n848, n849, n850, n851, n867, n868, n869, n870, n871, n872, n874,
         n875, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998;

  AOI21X1 U60 ( .A0(n123), .A1(n89), .B0(n90), .Y(n88) );
  AOI21X1 U72 ( .A0(n123), .A1(n98), .B0(n99), .Y(n97) );
  AOI21X1 U76 ( .A0(n114), .A1(n989), .B0(n103), .Y(n101) );
  AOI21X1 U88 ( .A0(n123), .A1(n988), .B0(n114), .Y(n110) );
  AOI21X1 U118 ( .A0(n160), .A1(n135), .B0(n136), .Y(n134) );
  AOI21X1 U132 ( .A0(n160), .A1(n313), .B0(n151), .Y(n145) );
  NOR2X2 U169 ( .A(n370), .B(n363), .Y(n170) );
  NOR2X2 U181 ( .A(n378), .B(n371), .Y(n183) );
  NOR2X2 U203 ( .A(n389), .B(n398), .Y(n199) );
  NOR2X2 U280 ( .A(n489), .B(n498), .Y(n248) );
  NAND2X4 U281 ( .A(n489), .B(n498), .Y(n249) );
  AOI21X1 U286 ( .A0(n961), .A1(n264), .B0(n259), .Y(n257) );
  ADDFHX4 U394 ( .A(n402), .B(n400), .CI(n391), .CO(n388), .S(n389) );
  ADDFHX4 U408 ( .A(n617), .B(n603), .CI(n432), .CO(n416), .S(n417) );
  ADDFHX4 U414 ( .A(n590), .B(n448), .CI(n446), .CO(n428), .S(n429) );
  ADDFHX4 U418 ( .A(n441), .B(n452), .CI(n439), .CO(n436), .S(n437) );
  ADDFHX4 U426 ( .A(n455), .B(n466), .CI(n453), .CO(n450), .S(n451) );
  ADDFHX4 U433 ( .A(n469), .B(n478), .CI(n467), .CO(n464), .S(n465) );
  ADDFHX4 U445 ( .A(n493), .B(n500), .CI(n491), .CO(n488), .S(n489) );
  OAI22X1 U478 ( .A0(n48), .A1(n693), .B0(n692), .B1(n46), .Y(n338) );
  OAI22X1 U479 ( .A0(n48), .A1(n694), .B0(n693), .B1(n46), .Y(n565) );
  OAI22X1 U480 ( .A0(n48), .A1(n695), .B0(n694), .B1(n46), .Y(n566) );
  OAI22X1 U481 ( .A0(n48), .A1(n696), .B0(n695), .B1(n46), .Y(n567) );
  OAI22X1 U483 ( .A0(n48), .A1(n698), .B0(n697), .B1(n46), .Y(n569) );
  OAI22X1 U485 ( .A0(n48), .A1(n700), .B0(n699), .B1(n46), .Y(n571) );
  OAI22X1 U488 ( .A0(n48), .A1(n703), .B0(n702), .B1(n46), .Y(n574) );
  OAI22X1 U492 ( .A0(n48), .A1(n707), .B0(n706), .B1(n46), .Y(n578) );
  OAI22X1 U528 ( .A0(n42), .A1(n724), .B0(n723), .B1(n40), .Y(n594) );
  OAI22X1 U547 ( .A0(n36), .A1(n870), .B0(n34), .B1(n742), .Y(n558) );
  OAI22X1 U550 ( .A0(n36), .A1(n727), .B0(n726), .B1(n34), .Y(n354) );
  OAI22X1 U551 ( .A0(n36), .A1(n728), .B0(n727), .B1(n34), .Y(n597) );
  OAI22X1 U552 ( .A0(n36), .A1(n729), .B0(n728), .B1(n34), .Y(n598) );
  OAI22X1 U554 ( .A0(n36), .A1(n731), .B0(n730), .B1(n34), .Y(n600) );
  OAI22X1 U555 ( .A0(n36), .A1(n732), .B0(n731), .B1(n34), .Y(n601) );
  OAI22X1 U556 ( .A0(n36), .A1(n733), .B0(n732), .B1(n34), .Y(n602) );
  OAI22X1 U557 ( .A0(n36), .A1(n734), .B0(n733), .B1(n34), .Y(n603) );
  OAI22X1 U558 ( .A0(n36), .A1(n735), .B0(n734), .B1(n34), .Y(n604) );
  OAI22X1 U559 ( .A0(n36), .A1(n736), .B0(n735), .B1(n34), .Y(n605) );
  OAI22X1 U562 ( .A0(n36), .A1(n739), .B0(n738), .B1(n34), .Y(n608) );
  OAI22X1 U563 ( .A0(n36), .A1(n740), .B0(n739), .B1(n34), .Y(n609) );
  OAI22X1 U564 ( .A0(n36), .A1(n741), .B0(n740), .B1(n34), .Y(n610) );
  OAI22X1 U583 ( .A0(n30), .A1(n871), .B0(n28), .B1(n759), .Y(n559) );
  OAI22X1 U586 ( .A0(n30), .A1(n744), .B0(n743), .B1(n28), .Y(n368) );
  OAI22X1 U587 ( .A0(n30), .A1(n745), .B0(n744), .B1(n28), .Y(n613) );
  OAI22X1 U588 ( .A0(n30), .A1(n746), .B0(n745), .B1(n28), .Y(n614) );
  OAI22X1 U589 ( .A0(n30), .A1(n747), .B0(n746), .B1(n28), .Y(n615) );
  OAI22X1 U590 ( .A0(n30), .A1(n748), .B0(n747), .B1(n28), .Y(n616) );
  OAI22X1 U591 ( .A0(n30), .A1(n749), .B0(n748), .B1(n28), .Y(n617) );
  OAI22X1 U592 ( .A0(n30), .A1(n750), .B0(n749), .B1(n28), .Y(n618) );
  OAI22X1 U593 ( .A0(n30), .A1(n751), .B0(n750), .B1(n28), .Y(n619) );
  OAI22X1 U594 ( .A0(n30), .A1(n752), .B0(n751), .B1(n28), .Y(n620) );
  OAI22X1 U595 ( .A0(n30), .A1(n753), .B0(n752), .B1(n28), .Y(n621) );
  OAI22X1 U596 ( .A0(n30), .A1(n754), .B0(n753), .B1(n28), .Y(n622) );
  OAI22X1 U597 ( .A0(n30), .A1(n755), .B0(n754), .B1(n28), .Y(n623) );
  OAI22X1 U599 ( .A0(n30), .A1(n757), .B0(n756), .B1(n28), .Y(n625) );
  OAI22X1 U600 ( .A0(n30), .A1(n758), .B0(n757), .B1(n28), .Y(n626) );
  OAI22X1 U658 ( .A0(n18), .A1(n778), .B0(n777), .B1(n16), .Y(n408) );
  OAI22X1 U662 ( .A0(n18), .A1(n782), .B0(n781), .B1(n16), .Y(n648) );
  OAI22X1 U664 ( .A0(n18), .A1(n784), .B0(n783), .B1(n16), .Y(n650) );
  OAI22X1 U668 ( .A0(n18), .A1(n788), .B0(n787), .B1(n16), .Y(n654) );
  OAI22X1 U670 ( .A0(n18), .A1(n790), .B0(n789), .B1(n16), .Y(n656) );
  OAI22X1 U691 ( .A0(n12), .A1(n874), .B0(n9), .B1(n810), .Y(n562) );
  OAI22X1 U696 ( .A0(n12), .A1(n797), .B0(n796), .B1(n9), .Y(n662) );
  OAI22X1 U698 ( .A0(n12), .A1(n799), .B0(n798), .B1(n9), .Y(n664) );
  OAI22X1 U700 ( .A0(n12), .A1(n801), .B0(n800), .B1(n9), .Y(n666) );
  OAI22X1 U701 ( .A0(n12), .A1(n802), .B0(n801), .B1(n9), .Y(n667) );
  OAI22X1 U702 ( .A0(n12), .A1(n803), .B0(n802), .B1(n9), .Y(n668) );
  OAI22X1 U703 ( .A0(n12), .A1(n804), .B0(n803), .B1(n9), .Y(n669) );
  OAI22X1 U704 ( .A0(n12), .A1(n805), .B0(n804), .B1(n9), .Y(n670) );
  OAI22X1 U705 ( .A0(n12), .A1(n806), .B0(n805), .B1(n9), .Y(n671) );
  OAI22X1 U706 ( .A0(n12), .A1(n807), .B0(n806), .B1(n9), .Y(n672) );
  OAI22X1 U707 ( .A0(n12), .A1(n808), .B0(n807), .B1(n9), .Y(n673) );
  OAI22X1 U708 ( .A0(n12), .A1(n809), .B0(n808), .B1(n9), .Y(n674) );
  OAI22X1 U731 ( .A0(n6), .A1(n813), .B0(n812), .B1(n867), .Y(n678) );
  OAI22X1 U732 ( .A0(n6), .A1(n814), .B0(n813), .B1(n867), .Y(n679) );
  OAI22X1 U733 ( .A0(n6), .A1(n815), .B0(n814), .B1(n867), .Y(n680) );
  OAI22X1 U735 ( .A0(n6), .A1(n817), .B0(n816), .B1(n867), .Y(n682) );
  OAI22X1 U737 ( .A0(n6), .A1(n819), .B0(n818), .B1(n867), .Y(n684) );
  OAI22X1 U739 ( .A0(n6), .A1(n821), .B0(n820), .B1(n867), .Y(n686) );
  OAI22X1 U740 ( .A0(n6), .A1(n822), .B0(n821), .B1(n867), .Y(n687) );
  OAI22X1 U741 ( .A0(n6), .A1(n823), .B0(n822), .B1(n867), .Y(n688) );
  OAI22X1 U742 ( .A0(n6), .A1(n824), .B0(n823), .B1(n867), .Y(n689) );
  OAI22X1 U743 ( .A0(n6), .A1(n825), .B0(n824), .B1(n867), .Y(n690) );
  OAI22X1 U744 ( .A0(n6), .A1(n826), .B0(n825), .B1(n867), .Y(n691) );
  NAND2X4 U786 ( .A(n46), .B(n844), .Y(n48) );
  XNOR2X4 U788 ( .A(n997), .B(a[14]), .Y(n46) );
  XNOR2X4 U791 ( .A(n996), .B(a[12]), .Y(n40) );
  NAND2X4 U792 ( .A(n34), .B(n846), .Y(n36) );
  XNOR2X4 U794 ( .A(n995), .B(a[10]), .Y(n34) );
  NAND2X4 U795 ( .A(n28), .B(n847), .Y(n30) );
  XNOR2X4 U797 ( .A(n994), .B(a[8]), .Y(n28) );
  NAND2X4 U798 ( .A(n22), .B(n848), .Y(n24) );
  NAND2X4 U801 ( .A(n16), .B(n849), .Y(n18) );
  XNOR2X4 U803 ( .A(n992), .B(a[4]), .Y(n16) );
  NAND2X4 U804 ( .A(n9), .B(n850), .Y(n12) );
  XNOR2X4 U806 ( .A(n991), .B(a[2]), .Y(n9) );
  NAND2X4 U807 ( .A(n851), .B(n867), .Y(n6) );
  ADDFHX4 U812 ( .A(n462), .B(n449), .CI(n460), .CO(n442), .S(n443) );
  AOI21X1 U813 ( .A0(n51), .A1(n193), .B0(n194), .Y(n192) );
  NOR2X4 U814 ( .A(n411), .B(n422), .Y(n211) );
  ADDFHX2 U815 ( .A(n427), .B(n438), .CI(n425), .CO(n422), .S(n423) );
  OAI22XL U816 ( .A0(n48), .A1(n868), .B0(n46), .B1(n708), .Y(n556) );
  XOR2X2 U817 ( .A(n201), .B(n64), .Y(product[20]) );
  BUFX20 U818 ( .A(a[3]), .Y(n992) );
  NAND2X4 U819 ( .A(n943), .B(n944), .Y(n945) );
  NAND2X4 U820 ( .A(n945), .B(n208), .Y(n51) );
  INVX2 U821 ( .A(n207), .Y(n943) );
  INVX1 U822 ( .A(n235), .Y(n944) );
  NAND2X1 U823 ( .A(n209), .B(n221), .Y(n207) );
  AOI21X2 U824 ( .A0(n255), .A1(n236), .B0(n237), .Y(n235) );
  AOI21X2 U825 ( .A0(n209), .A1(n222), .B0(n210), .Y(n208) );
  XOR2X2 U826 ( .A(n51), .B(n972), .Y(product[19]) );
  AOI21X1 U827 ( .A0(n51), .A1(n177), .B0(n178), .Y(n176) );
  AOI21X1 U828 ( .A0(n51), .A1(n168), .B0(n169), .Y(n167) );
  AOI21X1 U829 ( .A0(n51), .A1(n131), .B0(n132), .Y(n130) );
  AOI21X1 U830 ( .A0(n51), .A1(n142), .B0(n143), .Y(n141) );
  AOI21X1 U831 ( .A0(n51), .A1(n155), .B0(n156), .Y(n154) );
  AOI21X1 U832 ( .A0(n51), .A1(n186), .B0(n187), .Y(n185) );
  OR2X1 U833 ( .A(n12), .B(n800), .Y(n946) );
  OR2X1 U834 ( .A(n799), .B(n9), .Y(n947) );
  NAND2X2 U835 ( .A(n946), .B(n947), .Y(n665) );
  XNOR2XL U836 ( .A(b[9]), .B(n992), .Y(n800) );
  ADDFHX1 U837 ( .A(n637), .B(n665), .CI(n623), .CO(n494), .S(n495) );
  NOR2X2 U838 ( .A(n48), .B(n704), .Y(n948) );
  NOR2XL U839 ( .A(n703), .B(n46), .Y(n949) );
  OR2X4 U840 ( .A(n948), .B(n949), .Y(n575) );
  XNOR2XL U841 ( .A(b[4]), .B(n998), .Y(n703) );
  ADDFHX2 U842 ( .A(n575), .B(n434), .CI(n660), .CO(n420), .S(n421) );
  OR2X2 U843 ( .A(n30), .B(n756), .Y(n950) );
  OR2X1 U844 ( .A(n755), .B(n28), .Y(n951) );
  NAND2X4 U845 ( .A(n950), .B(n951), .Y(n624) );
  XNOR2XL U846 ( .A(b[2]), .B(n995), .Y(n756) );
  ADDFHX2 U847 ( .A(n638), .B(n624), .CI(n507), .CO(n502), .S(n503) );
  NAND2XL U848 ( .A(b[6]), .B(n993), .Y(n954) );
  NAND2X1 U849 ( .A(n952), .B(n953), .Y(n955) );
  NAND2X1 U850 ( .A(n954), .B(n955), .Y(n786) );
  CLKINVXL U851 ( .A(b[6]), .Y(n952) );
  CLKINVXL U852 ( .A(n993), .Y(n953) );
  BUFX12 U853 ( .A(a[5]), .Y(n993) );
  OAI22X1 U854 ( .A0(n24), .A1(n771), .B0(n770), .B1(n22), .Y(n638) );
  BUFX2 U855 ( .A(n607), .Y(n956) );
  OAI22X4 U856 ( .A0(n18), .A1(n786), .B0(n785), .B1(n16), .Y(n652) );
  OAI21XL U857 ( .A0(n254), .A1(n241), .B0(n242), .Y(n240) );
  OAI21X2 U858 ( .A0(n242), .A1(n238), .B0(n239), .Y(n237) );
  ADDFHX1 U859 ( .A(n622), .B(n594), .CI(n608), .CO(n482), .S(n483) );
  ADDFHX1 U860 ( .A(n604), .B(n646), .CI(n435), .CO(n432), .S(n433) );
  ADDHXL U861 ( .A(n681), .B(n652), .CO(n506), .S(n507) );
  ADDFHX1 U862 ( .A(n621), .B(n663), .CI(n649), .CO(n472), .S(n473) );
  ADDFHX1 U863 ( .A(n558), .B(n610), .CI(n666), .CO(n504), .S(n505) );
  AOI21X4 U864 ( .A0(n194), .A1(n181), .B0(n182), .Y(n52) );
  NOR2X2 U865 ( .A(n188), .B(n183), .Y(n181) );
  ADDFHX2 U866 ( .A(n415), .B(n424), .CI(n413), .CO(n410), .S(n411) );
  OAI22X1 U867 ( .A0(n12), .A1(n796), .B0(n795), .B1(n9), .Y(n661) );
  OR2XL U868 ( .A(n633), .B(n591), .Y(n448) );
  XNOR2X2 U869 ( .A(n633), .B(n591), .Y(n449) );
  ADDFHX1 U870 ( .A(n635), .B(n956), .CI(n486), .CO(n470), .S(n471) );
  OAI22XL U871 ( .A0(n36), .A1(n738), .B0(n737), .B1(n34), .Y(n607) );
  OAI22X2 U872 ( .A0(n42), .A1(n721), .B0(n720), .B1(n40), .Y(n591) );
  XNOR2X1 U873 ( .A(b[7]), .B(n993), .Y(n785) );
  XNOR2X1 U874 ( .A(b[7]), .B(n994), .Y(n768) );
  XNOR2X1 U875 ( .A(b[4]), .B(n997), .Y(n720) );
  OAI22X2 U876 ( .A0(n12), .A1(n795), .B0(n794), .B1(n9), .Y(n434) );
  BUFX2 U877 ( .A(n661), .Y(n957) );
  ADDFHX1 U878 ( .A(n602), .B(n630), .CI(n409), .CO(n406), .S(n407) );
  XNOR2X1 U879 ( .A(b[2]), .B(n996), .Y(n739) );
  XNOR2X1 U880 ( .A(b[2]), .B(n997), .Y(n722) );
  INVX1 U881 ( .A(n434), .Y(n435) );
  ADDFHX1 U882 ( .A(n662), .B(n606), .CI(n620), .CO(n458), .S(n459) );
  OAI22X2 U883 ( .A0(n24), .A1(n766), .B0(n765), .B1(n22), .Y(n633) );
  NAND2X4 U884 ( .A(n40), .B(n845), .Y(n42) );
  XOR2X2 U885 ( .A(n997), .B(a[12]), .Y(n845) );
  ADDFHX1 U886 ( .A(n619), .B(n957), .CI(n676), .CO(n446), .S(n447) );
  AOI21XL U887 ( .A0(n51), .A1(n94), .B0(n95), .Y(n93) );
  AOI21XL U888 ( .A0(n51), .A1(n118), .B0(n119), .Y(n117) );
  AOI21XL U889 ( .A0(n51), .A1(n107), .B0(n108), .Y(n106) );
  AOI21XL U890 ( .A0(n51), .A1(n319), .B0(n203), .Y(n201) );
  XNOR2X2 U891 ( .A(b[11]), .B(n992), .Y(n798) );
  XNOR2X1 U892 ( .A(b[11]), .B(n993), .Y(n781) );
  OAI21X4 U893 ( .A0(n227), .A1(n233), .B0(n228), .Y(n222) );
  NOR2X4 U894 ( .A(n437), .B(n450), .Y(n227) );
  XNOR2X2 U895 ( .A(b[8]), .B(n994), .Y(n767) );
  XNOR2X1 U896 ( .A(b[8]), .B(n993), .Y(n784) );
  XNOR2X1 U897 ( .A(b[8]), .B(n991), .Y(n818) );
  XNOR2X2 U898 ( .A(b[12]), .B(n992), .Y(n797) );
  XNOR2X2 U899 ( .A(b[12]), .B(n991), .Y(n814) );
  XNOR2X1 U900 ( .A(b[12]), .B(n993), .Y(n780) );
  XNOR2X2 U901 ( .A(b[12]), .B(n994), .Y(n763) );
  XNOR2X2 U902 ( .A(b[9]), .B(n994), .Y(n766) );
  XNOR2X1 U903 ( .A(b[9]), .B(n993), .Y(n783) );
  XNOR2X2 U904 ( .A(b[9]), .B(n991), .Y(n817) );
  XNOR2X1 U905 ( .A(b[9]), .B(n996), .Y(n732) );
  XNOR2X2 U906 ( .A(b[15]), .B(n991), .Y(n811) );
  XNOR2X1 U907 ( .A(b[15]), .B(n992), .Y(n794) );
  XNOR2X1 U908 ( .A(b[15]), .B(n993), .Y(n777) );
  XNOR2X2 U909 ( .A(b[13]), .B(n992), .Y(n796) );
  XNOR2X2 U910 ( .A(b[13]), .B(n991), .Y(n813) );
  XNOR2X1 U911 ( .A(b[13]), .B(n993), .Y(n779) );
  XNOR2X2 U912 ( .A(b[13]), .B(n994), .Y(n762) );
  XNOR2X2 U913 ( .A(b[14]), .B(n992), .Y(n795) );
  XNOR2X2 U914 ( .A(b[14]), .B(n991), .Y(n812) );
  BUFX8 U915 ( .A(a[9]), .Y(n995) );
  BUFX8 U916 ( .A(a[11]), .Y(n996) );
  BUFX8 U917 ( .A(a[13]), .Y(n997) );
  XOR2X1 U918 ( .A(n994), .B(a[6]), .Y(n848) );
  ADDFX2 U919 ( .A(n584), .B(n570), .CI(n369), .CO(n366), .S(n367) );
  ADDFX2 U920 ( .A(n354), .B(n567), .CI(n596), .CO(n348), .S(n349) );
  ADDFX2 U921 ( .A(n582), .B(n568), .CI(n355), .CO(n352), .S(n353) );
  ADDFHX1 U922 ( .A(n392), .B(n390), .CI(n381), .CO(n378), .S(n379) );
  ADDFHX1 U923 ( .A(n367), .B(n365), .CI(n372), .CO(n362), .S(n363) );
  ADDFHX1 U924 ( .A(n382), .B(n373), .CI(n380), .CO(n370), .S(n371) );
  NAND2X2 U925 ( .A(n399), .B(n410), .Y(n205) );
  NOR2X1 U926 ( .A(n379), .B(n388), .Y(n188) );
  OAI21X1 U927 ( .A0(n158), .A1(n124), .B0(n125), .Y(n123) );
  ADDHXL U928 ( .A(n687), .B(n658), .CO(n542), .S(n543) );
  ADDFHX1 U929 ( .A(n557), .B(n664), .CI(n636), .CO(n484), .S(n485) );
  OAI22X1 U930 ( .A0(n42), .A1(n869), .B0(n40), .B1(n725), .Y(n557) );
  XNOR2X1 U931 ( .A(n81), .B(n303), .Y(product[3]) );
  ADDFHX1 U932 ( .A(n513), .B(n518), .CI(n511), .CO(n508), .S(n509) );
  ADDFHX1 U933 ( .A(n503), .B(n510), .CI(n501), .CO(n498), .S(n499) );
  NAND2X1 U934 ( .A(n509), .B(n516), .Y(n266) );
  ADDFHX1 U935 ( .A(n556), .B(n578), .CI(n592), .CO(n460), .S(n461) );
  ADDFX2 U936 ( .A(n585), .B(n599), .CI(n613), .CO(n374), .S(n375) );
  ADDFX1 U937 ( .A(n573), .B(n408), .CI(n644), .CO(n396), .S(n397) );
  ADDFX2 U938 ( .A(n586), .B(n614), .CI(n387), .CO(n384), .S(n385) );
  ADDFX2 U939 ( .A(n629), .B(n587), .CI(n601), .CO(n394), .S(n395) );
  BUFX8 U940 ( .A(a[15]), .Y(n998) );
  NOR2X1 U941 ( .A(n271), .B(n274), .Y(n269) );
  OAI21XL U942 ( .A0(n271), .A1(n275), .B0(n272), .Y(n270) );
  INVX2 U943 ( .A(n266), .Y(n264) );
  ADDFX2 U944 ( .A(n597), .B(n583), .CI(n366), .CO(n358), .S(n359) );
  NOR2X1 U945 ( .A(n399), .B(n410), .Y(n204) );
  NAND2X2 U946 ( .A(n451), .B(n464), .Y(n233) );
  NOR2X1 U947 ( .A(n356), .B(n351), .Y(n148) );
  ADDFX2 U948 ( .A(n361), .B(n359), .CI(n364), .CO(n356), .S(n357) );
  ADDFX2 U949 ( .A(n360), .B(n353), .CI(n358), .CO(n350), .S(n351) );
  NAND2X1 U950 ( .A(n159), .B(n135), .Y(n133) );
  ADDFX2 U951 ( .A(n581), .B(n352), .CI(n349), .CO(n346), .S(n347) );
  NAND2X1 U952 ( .A(n122), .B(n98), .Y(n96) );
  NOR2X1 U953 ( .A(n204), .B(n199), .Y(n193) );
  NOR2X1 U954 ( .A(n157), .B(n124), .Y(n122) );
  NAND2X1 U955 ( .A(n356), .B(n351), .Y(n149) );
  INVX2 U956 ( .A(n166), .Y(n164) );
  NOR2BXL U957 ( .AN(n193), .B(n188), .Y(n186) );
  NAND2X1 U958 ( .A(n370), .B(n363), .Y(n171) );
  CLKINVXL U959 ( .A(n53), .Y(n177) );
  NOR2X1 U960 ( .A(n350), .B(n347), .Y(n137) );
  NOR2X1 U961 ( .A(n346), .B(n343), .Y(n128) );
  BUFX8 U962 ( .A(n52), .Y(n990) );
  ADDHXL U963 ( .A(n689), .B(n562), .CO(n546), .S(n547) );
  ADDFX2 U964 ( .A(n643), .B(n686), .CI(n657), .CO(n538), .S(n539) );
  ADDHXL U965 ( .A(n685), .B(n656), .CO(n534), .S(n535) );
  ADDFX2 U966 ( .A(n611), .B(n682), .CI(n625), .CO(n514), .S(n515) );
  NAND2X1 U967 ( .A(n547), .B(n674), .Y(n302) );
  OAI21X1 U968 ( .A0(n304), .A1(n307), .B0(n305), .Y(n303) );
  ADDFX2 U969 ( .A(n561), .B(n672), .CI(n543), .CO(n540), .S(n541) );
  OR2X1 U970 ( .A(n541), .B(n544), .Y(n987) );
  ADDFX2 U971 ( .A(n529), .B(n532), .CI(n527), .CO(n524), .S(n525) );
  ADDFX2 U972 ( .A(n559), .B(n626), .CI(n640), .CO(n520), .S(n521) );
  ADDFX2 U973 ( .A(n668), .B(n523), .CI(n528), .CO(n518), .S(n519) );
  ADDFHX1 U974 ( .A(n522), .B(n515), .CI(n520), .CO(n510), .S(n511) );
  NAND2BX1 U975 ( .AN(b[0]), .B(n998), .Y(n708) );
  ADDFX2 U976 ( .A(n651), .B(n506), .CI(n497), .CO(n492), .S(n493) );
  NAND2X1 U977 ( .A(n691), .B(n563), .Y(n307) );
  ADDFX2 U978 ( .A(n504), .B(n502), .CI(n495), .CO(n490), .S(n491) );
  ADDFX2 U979 ( .A(n487), .B(n496), .CI(n494), .CO(n480), .S(n481) );
  NOR2X1 U980 ( .A(n517), .B(n524), .Y(n271) );
  NOR2X1 U981 ( .A(n525), .B(n530), .Y(n274) );
  NAND2X1 U982 ( .A(n525), .B(n530), .Y(n275) );
  ADDFX2 U983 ( .A(n634), .B(n463), .CI(n474), .CO(n456), .S(n457) );
  ADDFX2 U984 ( .A(n475), .B(n484), .CI(n473), .CO(n468), .S(n469) );
  ADDFX2 U985 ( .A(n485), .B(n483), .CI(n492), .CO(n478), .S(n479) );
  ADDFX2 U986 ( .A(n472), .B(n470), .CI(n459), .CO(n454), .S(n455) );
  ADDFX2 U987 ( .A(n482), .B(n471), .CI(n480), .CO(n466), .S(n467) );
  ADDFX2 U988 ( .A(n418), .B(n416), .CI(n414), .CO(n400), .S(n401) );
  ADDFX2 U989 ( .A(n420), .B(n405), .CI(n407), .CO(n402), .S(n403) );
  ADDFHX1 U990 ( .A(n481), .B(n490), .CI(n479), .CO(n476), .S(n477) );
  ADDFX2 U991 ( .A(n430), .B(n421), .CI(n419), .CO(n414), .S(n415) );
  ADDFX2 U992 ( .A(n428), .B(n417), .CI(n426), .CO(n412), .S(n413) );
  ADDFX2 U993 ( .A(n461), .B(n457), .CI(n468), .CO(n452), .S(n453) );
  ADDFX2 U994 ( .A(n458), .B(n447), .CI(n445), .CO(n440), .S(n441) );
  ADDFHX1 U995 ( .A(n456), .B(n443), .CI(n454), .CO(n438), .S(n439) );
  ADDFHX1 U996 ( .A(n444), .B(n433), .CI(n431), .CO(n426), .S(n427) );
  ADDFX2 U997 ( .A(n442), .B(n429), .CI(n440), .CO(n424), .S(n425) );
  XNOR2X1 U998 ( .A(n247), .B(n71), .Y(product[13]) );
  OAI21X1 U999 ( .A0(n254), .A1(n248), .B0(n249), .Y(n247) );
  ADDFX2 U1000 ( .A(n615), .B(n406), .CI(n404), .CO(n392), .S(n393) );
  ADDFX2 U1001 ( .A(n395), .B(n397), .CI(n393), .CO(n390), .S(n391) );
  ADDFX2 U1002 ( .A(n598), .B(n376), .CI(n374), .CO(n364), .S(n365) );
  ADDFX2 U1003 ( .A(n384), .B(n377), .CI(n375), .CO(n372), .S(n373) );
  ADDFX2 U1004 ( .A(n394), .B(n385), .CI(n383), .CO(n380), .S(n381) );
  ADDFHX1 U1005 ( .A(n403), .B(n412), .CI(n401), .CO(n398), .S(n399) );
  XOR2X1 U1006 ( .A(a[14]), .B(n998), .Y(n844) );
  NOR2X1 U1007 ( .A(n137), .B(n128), .Y(n126) );
  NAND2X1 U1008 ( .A(n313), .B(n126), .Y(n124) );
  NOR2X2 U1009 ( .A(n465), .B(n476), .Y(n238) );
  AOI21X2 U1010 ( .A0(n960), .A1(n251), .B0(n244), .Y(n242) );
  INVX2 U1011 ( .A(n249), .Y(n251) );
  NAND2X1 U1012 ( .A(n960), .B(n326), .Y(n241) );
  NAND2X1 U1013 ( .A(n465), .B(n476), .Y(n239) );
  NAND2X1 U1014 ( .A(n961), .B(n983), .Y(n256) );
  INVX2 U1015 ( .A(a[0]), .Y(n867) );
  XOR2X1 U1016 ( .A(n213), .B(n66), .Y(product[18]) );
  NAND2X1 U1017 ( .A(n320), .B(n212), .Y(n66) );
  XOR2X1 U1018 ( .A(n229), .B(n68), .Y(product[16]) );
  XOR2X1 U1019 ( .A(n220), .B(n67), .Y(product[17]) );
  NAND2X1 U1020 ( .A(n321), .B(n219), .Y(n67) );
  INVX2 U1021 ( .A(n158), .Y(n160) );
  NAND2X1 U1022 ( .A(n411), .B(n422), .Y(n212) );
  NAND2X1 U1023 ( .A(n423), .B(n436), .Y(n219) );
  NOR2X1 U1024 ( .A(n227), .B(n232), .Y(n221) );
  NOR2X1 U1025 ( .A(n53), .B(n120), .Y(n118) );
  AND2X1 U1026 ( .A(n319), .B(n205), .Y(n972) );
  XOR2X1 U1027 ( .A(n192), .B(n63), .Y(product[21]) );
  XOR2X1 U1028 ( .A(n154), .B(n59), .Y(product[25]) );
  OAI21X1 U1029 ( .A0(n990), .A1(n157), .B0(n158), .Y(n156) );
  XOR2X1 U1030 ( .A(n167), .B(n60), .Y(product[24]) );
  NOR2X1 U1031 ( .A(n53), .B(n109), .Y(n107) );
  XOR2X1 U1032 ( .A(n185), .B(n62), .Y(product[22]) );
  XOR2X1 U1033 ( .A(n176), .B(n973), .Y(product[23]) );
  XNOR2X1 U1034 ( .A(n141), .B(n975), .Y(product[26]) );
  XNOR2X1 U1035 ( .A(n130), .B(n976), .Y(product[27]) );
  XNOR2X1 U1036 ( .A(n93), .B(n981), .Y(product[30]) );
  INVX2 U1037 ( .A(n91), .Y(n308) );
  NOR2X1 U1038 ( .A(n53), .B(n87), .Y(n85) );
  XNOR2X1 U1039 ( .A(n240), .B(n70), .Y(product[14]) );
  BUFX2 U1040 ( .A(n653), .Y(n958) );
  AND2X2 U1041 ( .A(n984), .B(n986), .Y(n959) );
  OR2X2 U1042 ( .A(n477), .B(n488), .Y(n960) );
  AOI21X1 U1043 ( .A0(n295), .A1(n987), .B0(n292), .Y(n290) );
  OR2X1 U1044 ( .A(n499), .B(n508), .Y(n961) );
  AND2X1 U1045 ( .A(n978), .B(n307), .Y(product[1]) );
  AOI21XL U1046 ( .A0(n51), .A1(n85), .B0(n86), .Y(product[31]) );
  OAI22X1 U1047 ( .A0(n18), .A1(n792), .B0(n791), .B1(n16), .Y(n658) );
  NAND2X1 U1048 ( .A(n993), .B(a[6]), .Y(n965) );
  NAND2X2 U1049 ( .A(n963), .B(n964), .Y(n966) );
  NAND2X4 U1050 ( .A(n965), .B(n966), .Y(n22) );
  INVX2 U1051 ( .A(n993), .Y(n963) );
  INVX2 U1052 ( .A(a[6]), .Y(n964) );
  NOR2BX1 U1053 ( .AN(b[0]), .B(n22), .Y(n643) );
  OAI22XL U1054 ( .A0(n24), .A1(n774), .B0(n773), .B1(n22), .Y(n641) );
  OAI22XL U1055 ( .A0(n24), .A1(n768), .B0(n767), .B1(n22), .Y(n635) );
  OAI22XL U1056 ( .A0(n24), .A1(n769), .B0(n768), .B1(n22), .Y(n636) );
  OAI22XL U1057 ( .A0(n24), .A1(n767), .B0(n766), .B1(n22), .Y(n634) );
  OAI22XL U1058 ( .A0(n24), .A1(n764), .B0(n763), .B1(n22), .Y(n631) );
  OAI22X1 U1059 ( .A0(n24), .A1(n872), .B0(n22), .B1(n776), .Y(n560) );
  OAI22XL U1060 ( .A0(n24), .A1(n772), .B0(n771), .B1(n22), .Y(n639) );
  OAI22XL U1061 ( .A0(n24), .A1(n770), .B0(n769), .B1(n22), .Y(n637) );
  OAI22XL U1062 ( .A0(n24), .A1(n773), .B0(n772), .B1(n22), .Y(n640) );
  OAI22XL U1063 ( .A0(n24), .A1(n765), .B0(n764), .B1(n22), .Y(n632) );
  OAI22XL U1064 ( .A0(n24), .A1(n761), .B0(n760), .B1(n22), .Y(n386) );
  OAI22XL U1065 ( .A0(n24), .A1(n762), .B0(n761), .B1(n22), .Y(n629) );
  NAND2X2 U1066 ( .A(n959), .B(n967), .Y(n968) );
  NAND2X2 U1067 ( .A(n968), .B(n279), .Y(n277) );
  CLKINVX2 U1068 ( .A(n290), .Y(n967) );
  INVX1 U1069 ( .A(n277), .Y(n276) );
  OR2X1 U1070 ( .A(n547), .B(n674), .Y(n985) );
  XNOR2XL U1071 ( .A(b[1]), .B(n994), .Y(n774) );
  CLKINVXL U1072 ( .A(n990), .Y(n178) );
  NAND2X1 U1073 ( .A(n159), .B(n313), .Y(n144) );
  NAND2BX1 U1074 ( .AN(b[0]), .B(n996), .Y(n742) );
  INVX3 U1075 ( .A(n255), .Y(n254) );
  INVX1 U1076 ( .A(n232), .Y(n323) );
  NOR2XL U1077 ( .A(n24), .B(n775), .Y(n969) );
  NOR2XL U1078 ( .A(n774), .B(n22), .Y(n970) );
  OR2X1 U1079 ( .A(n969), .B(n970), .Y(n642) );
  XNOR2XL U1080 ( .A(b[0]), .B(n994), .Y(n775) );
  NOR2X1 U1081 ( .A(n53), .B(n170), .Y(n168) );
  XOR2X1 U1082 ( .A(n996), .B(a[10]), .Y(n846) );
  OAI21X2 U1083 ( .A0(n211), .A1(n219), .B0(n212), .Y(n210) );
  NAND2BX1 U1084 ( .AN(n199), .B(n200), .Y(n64) );
  OAI21X2 U1085 ( .A0(n199), .A1(n205), .B0(n200), .Y(n194) );
  INVX1 U1086 ( .A(n261), .Y(n259) );
  NAND2X1 U1087 ( .A(n315), .B(n982), .Y(n157) );
  NAND2X1 U1088 ( .A(n517), .B(n524), .Y(n272) );
  AOI21X1 U1089 ( .A0(n985), .A1(n303), .B0(n300), .Y(n298) );
  OR2XL U1090 ( .A(n691), .B(n563), .Y(n978) );
  AOI21X1 U1091 ( .A0(n214), .A1(n234), .B0(n215), .Y(n213) );
  XOR2X1 U1092 ( .A(n234), .B(n971), .Y(product[15]) );
  AND2X1 U1093 ( .A(n323), .B(n233), .Y(n971) );
  AOI21XL U1094 ( .A0(n234), .A1(n323), .B0(n231), .Y(n229) );
  NAND2XL U1095 ( .A(n324), .B(n239), .Y(n70) );
  AOI21X2 U1096 ( .A0(n269), .A1(n277), .B0(n270), .Y(n268) );
  AOI21X1 U1097 ( .A0(n267), .A1(n983), .B0(n264), .Y(n262) );
  NAND2X2 U1098 ( .A(n437), .B(n450), .Y(n228) );
  INVX1 U1099 ( .A(n170), .Y(n315) );
  CLKINVXL U1100 ( .A(n982), .Y(n979) );
  INVX2 U1101 ( .A(n148), .Y(n313) );
  INVX1 U1102 ( .A(n283), .Y(n281) );
  NAND2X1 U1103 ( .A(n477), .B(n488), .Y(n246) );
  OR2XL U1104 ( .A(n537), .B(n540), .Y(n986) );
  NAND2XL U1105 ( .A(n541), .B(n544), .Y(n294) );
  XNOR2XL U1106 ( .A(b[0]), .B(n991), .Y(n826) );
  XOR2X2 U1107 ( .A(n991), .B(a[0]), .Y(n851) );
  XNOR2XL U1108 ( .A(b[3]), .B(n997), .Y(n721) );
  XNOR2XL U1109 ( .A(b[3]), .B(n998), .Y(n704) );
  XNOR2XL U1110 ( .A(b[7]), .B(n997), .Y(n717) );
  XNOR2XL U1111 ( .A(b[8]), .B(n997), .Y(n716) );
  XNOR2XL U1112 ( .A(b[9]), .B(n997), .Y(n715) );
  XNOR2XL U1113 ( .A(b[10]), .B(n997), .Y(n714) );
  XNOR2XL U1114 ( .A(b[11]), .B(n998), .Y(n696) );
  XNOR2XL U1115 ( .A(b[12]), .B(n998), .Y(n695) );
  NOR2XL U1116 ( .A(n53), .B(n144), .Y(n142) );
  NOR2XL U1117 ( .A(n53), .B(n96), .Y(n94) );
  NAND2BX1 U1118 ( .AN(n227), .B(n228), .Y(n68) );
  AOI21XL U1119 ( .A0(n234), .A1(n221), .B0(n222), .Y(n220) );
  XOR2X1 U1120 ( .A(n254), .B(n72), .Y(product[12]) );
  XOR2X1 U1121 ( .A(n262), .B(n73), .Y(product[11]) );
  XNOR2X1 U1122 ( .A(n273), .B(n75), .Y(product[9]) );
  NAND2X1 U1123 ( .A(n329), .B(n272), .Y(n75) );
  OAI21XL U1124 ( .A0(n276), .A1(n274), .B0(n275), .Y(n273) );
  XOR2X1 U1125 ( .A(n276), .B(n76), .Y(product[8]) );
  NAND2XL U1126 ( .A(n330), .B(n275), .Y(n76) );
  NAND2XL U1127 ( .A(n316), .B(n184), .Y(n62) );
  NAND2BXL U1128 ( .AN(n188), .B(n191), .Y(n63) );
  NAND2XL U1129 ( .A(n315), .B(n171), .Y(n973) );
  NAND2X1 U1130 ( .A(n389), .B(n398), .Y(n200) );
  INVX2 U1131 ( .A(n149), .Y(n151) );
  NAND2XL U1132 ( .A(n122), .B(n89), .Y(n87) );
  NAND2XL U1133 ( .A(n499), .B(n508), .Y(n261) );
  XOR2X1 U1134 ( .A(n974), .B(n967), .Y(product[6]) );
  AND2X1 U1135 ( .A(n986), .B(n288), .Y(n974) );
  XOR2X1 U1136 ( .A(n284), .B(n77), .Y(product[7]) );
  AOI21XL U1137 ( .A0(n967), .A1(n986), .B0(n286), .Y(n284) );
  XOR2XL U1138 ( .A(n80), .B(n298), .Y(product[4]) );
  CLKINVXL U1139 ( .A(n296), .Y(n334) );
  XNOR2XL U1140 ( .A(n79), .B(n295), .Y(product[5]) );
  NAND2XL U1141 ( .A(n987), .B(n294), .Y(n79) );
  AND2X1 U1142 ( .A(n312), .B(n140), .Y(n975) );
  XOR2XL U1143 ( .A(n82), .B(n307), .Y(product[2]) );
  NAND2XL U1144 ( .A(n336), .B(n305), .Y(n82) );
  CLKINVXL U1145 ( .A(n304), .Y(n336) );
  AND2X1 U1146 ( .A(n311), .B(n129), .Y(n976) );
  AOI21XL U1147 ( .A0(n126), .A1(n151), .B0(n127), .Y(n125) );
  XOR2X1 U1148 ( .A(n106), .B(n977), .Y(product[29]) );
  NAND2X1 U1149 ( .A(n989), .B(n105), .Y(n977) );
  NAND2X1 U1150 ( .A(n122), .B(n988), .Y(n109) );
  XOR2X1 U1151 ( .A(n117), .B(n56), .Y(product[28]) );
  NAND2XL U1152 ( .A(n362), .B(n357), .Y(n166) );
  NOR2X1 U1153 ( .A(n148), .B(n137), .Y(n135) );
  ADDFHX1 U1154 ( .A(n514), .B(n512), .CI(n505), .CO(n500), .S(n501) );
  OR2X2 U1155 ( .A(n531), .B(n536), .Y(n984) );
  NAND2XL U1156 ( .A(n531), .B(n536), .Y(n283) );
  ADDFHX2 U1157 ( .A(n521), .B(n526), .CI(n519), .CO(n516), .S(n517) );
  NAND2XL U1158 ( .A(n537), .B(n540), .Y(n288) );
  NAND2XL U1159 ( .A(n545), .B(n546), .Y(n297) );
  NAND2XL U1160 ( .A(n350), .B(n347), .Y(n140) );
  OAI22X1 U1161 ( .A0(n6), .A1(n875), .B0(n827), .B1(n867), .Y(n563) );
  CLKINVXL U1162 ( .A(n991), .Y(n875) );
  CLKINVXL U1163 ( .A(n992), .Y(n874) );
  OAI22XL U1164 ( .A0(n6), .A1(n820), .B0(n819), .B1(n867), .Y(n685) );
  OAI22XL U1165 ( .A0(n18), .A1(n963), .B0(n16), .B1(n793), .Y(n561) );
  OAI22XL U1166 ( .A0(n6), .A1(n816), .B0(n815), .B1(n867), .Y(n681) );
  NAND2BXL U1167 ( .AN(b[0]), .B(n994), .Y(n776) );
  NAND2BXL U1168 ( .AN(b[0]), .B(n992), .Y(n810) );
  OAI22XL U1169 ( .A0(n36), .A1(n737), .B0(n736), .B1(n34), .Y(n606) );
  OAI22XL U1170 ( .A0(n12), .A1(n798), .B0(n797), .B1(n9), .Y(n663) );
  OAI22XL U1171 ( .A0(n48), .A1(n706), .B0(n705), .B1(n46), .Y(n577) );
  OAI22XL U1172 ( .A0(n18), .A1(n780), .B0(n779), .B1(n16), .Y(n646) );
  CLKINVXL U1173 ( .A(n994), .Y(n872) );
  ADDHX1 U1174 ( .A(n677), .B(n648), .CO(n462), .S(n463) );
  OAI22XL U1175 ( .A0(n6), .A1(n812), .B0(n811), .B1(n867), .Y(n677) );
  CLKINVXL U1176 ( .A(n996), .Y(n870) );
  CLKINVXL U1177 ( .A(n995), .Y(n871) );
  OAI22XL U1178 ( .A0(n48), .A1(n705), .B0(n704), .B1(n46), .Y(n576) );
  INVX1 U1179 ( .A(n408), .Y(n409) );
  OAI22XL U1180 ( .A0(n24), .A1(n763), .B0(n762), .B1(n22), .Y(n630) );
  CLKINVXL U1181 ( .A(n794), .Y(n554) );
  CLKINVXL U1182 ( .A(n760), .Y(n552) );
  CLKINVXL U1183 ( .A(n777), .Y(n553) );
  OAI22XL U1184 ( .A0(n48), .A1(n702), .B0(n701), .B1(n46), .Y(n573) );
  ADDFHX2 U1185 ( .A(n600), .B(n572), .CI(n396), .CO(n382), .S(n383) );
  OAI22XL U1186 ( .A0(n48), .A1(n701), .B0(n700), .B1(n46), .Y(n572) );
  INVXL U1187 ( .A(n368), .Y(n369) );
  OAI22XL U1188 ( .A0(n48), .A1(n699), .B0(n698), .B1(n46), .Y(n570) );
  OAI22XL U1189 ( .A0(n36), .A1(n730), .B0(n729), .B1(n34), .Y(n599) );
  CLKINVXL U1190 ( .A(n997), .Y(n869) );
  CLKINVXL U1191 ( .A(n998), .Y(n868) );
  OAI22XL U1192 ( .A0(n48), .A1(n697), .B0(n696), .B1(n46), .Y(n568) );
  XNOR2X1 U1193 ( .A(b[1]), .B(n997), .Y(n723) );
  XNOR2X1 U1194 ( .A(b[1]), .B(n998), .Y(n706) );
  XNOR2X1 U1195 ( .A(b[2]), .B(n998), .Y(n705) );
  XNOR2X1 U1196 ( .A(b[6]), .B(n997), .Y(n718) );
  XNOR2X1 U1197 ( .A(b[5]), .B(n997), .Y(n719) );
  XNOR2X1 U1198 ( .A(b[5]), .B(n998), .Y(n702) );
  XNOR2X1 U1199 ( .A(b[6]), .B(n998), .Y(n701) );
  XNOR2X1 U1200 ( .A(b[8]), .B(n998), .Y(n699) );
  XNOR2X1 U1201 ( .A(b[7]), .B(n998), .Y(n700) );
  XNOR2X1 U1202 ( .A(b[9]), .B(n998), .Y(n698) );
  XNOR2XL U1203 ( .A(b[15]), .B(n995), .Y(n743) );
  XNOR2X1 U1204 ( .A(b[10]), .B(n998), .Y(n697) );
  INVX2 U1205 ( .A(n235), .Y(n234) );
  INVX2 U1206 ( .A(n122), .Y(n120) );
  CLKINVXL U1207 ( .A(n211), .Y(n320) );
  CLKINVXL U1208 ( .A(n216), .Y(n321) );
  NAND2X2 U1209 ( .A(n193), .B(n181), .Y(n53) );
  INVX2 U1210 ( .A(n268), .Y(n267) );
  CLKINVXL U1211 ( .A(n222), .Y(n224) );
  OAI21XL U1212 ( .A0(n990), .A1(n144), .B0(n145), .Y(n143) );
  NOR2XL U1213 ( .A(n53), .B(n133), .Y(n131) );
  NOR2BXL U1214 ( .AN(n221), .B(n216), .Y(n214) );
  INVX2 U1215 ( .A(n157), .Y(n159) );
  CLKINVXL U1216 ( .A(n233), .Y(n231) );
  CLKINVXL U1217 ( .A(n204), .Y(n319) );
  CLKINVXL U1218 ( .A(n205), .Y(n203) );
  AOI2BB1X4 U1219 ( .A0N(n979), .A1N(n171), .B0(n164), .Y(n158) );
  OAI21XL U1220 ( .A0(n990), .A1(n96), .B0(n97), .Y(n95) );
  INVX2 U1221 ( .A(n101), .Y(n99) );
  OAI21XL U1222 ( .A0(n990), .A1(n87), .B0(n88), .Y(n86) );
  INVX2 U1223 ( .A(n246), .Y(n244) );
  CLKINVXL U1224 ( .A(n183), .Y(n316) );
  INVX2 U1225 ( .A(n248), .Y(n326) );
  OAI21X1 U1226 ( .A0(n183), .A1(n191), .B0(n184), .Y(n182) );
  NAND2X1 U1227 ( .A(n313), .B(n149), .Y(n59) );
  NOR2XL U1228 ( .A(n53), .B(n157), .Y(n155) );
  NAND2XL U1229 ( .A(n960), .B(n246), .Y(n71) );
  CLKINVXL U1230 ( .A(n271), .Y(n329) );
  NAND2XL U1231 ( .A(n961), .B(n261), .Y(n73) );
  OAI21XL U1232 ( .A0(n990), .A1(n170), .B0(n171), .Y(n169) );
  NAND2X1 U1233 ( .A(n982), .B(n166), .Y(n60) );
  NOR2X2 U1234 ( .A(n451), .B(n464), .Y(n232) );
  NAND2XL U1235 ( .A(n326), .B(n249), .Y(n72) );
  OAI21XL U1236 ( .A0(n990), .A1(n120), .B0(n121), .Y(n119) );
  CLKINVXL U1237 ( .A(n123), .Y(n121) );
  CLKINVXL U1238 ( .A(n274), .Y(n330) );
  OAI21XL U1239 ( .A0(n196), .A1(n188), .B0(n191), .Y(n187) );
  CLKINVXL U1240 ( .A(n194), .Y(n196) );
  XOR2X1 U1241 ( .A(n267), .B(n980), .Y(product[10]) );
  AND2X1 U1242 ( .A(n983), .B(n266), .Y(n980) );
  INVX2 U1243 ( .A(n100), .Y(n98) );
  OAI21XL U1244 ( .A0(n140), .A1(n128), .B0(n129), .Y(n127) );
  AND2X1 U1245 ( .A(n308), .B(n92), .Y(n981) );
  OR2X4 U1246 ( .A(n362), .B(n357), .Y(n982) );
  OAI21XL U1247 ( .A0(n990), .A1(n109), .B0(n110), .Y(n108) );
  OAI21X1 U1248 ( .A0(n101), .A1(n91), .B0(n92), .Y(n90) );
  AOI21X1 U1249 ( .A0(n984), .A1(n286), .B0(n281), .Y(n279) );
  CLKINVXL U1250 ( .A(n128), .Y(n311) );
  OAI21XL U1251 ( .A0(n990), .A1(n133), .B0(n134), .Y(n132) );
  OAI21XL U1252 ( .A0(n149), .A1(n137), .B0(n140), .Y(n136) );
  NAND2X1 U1253 ( .A(n988), .B(n116), .Y(n56) );
  INVX2 U1254 ( .A(n302), .Y(n300) );
  OAI21X1 U1255 ( .A0(n298), .A1(n296), .B0(n297), .Y(n295) );
  INVX2 U1256 ( .A(n294), .Y(n292) );
  NAND2X1 U1257 ( .A(n985), .B(n302), .Y(n81) );
  CLKINVXL U1258 ( .A(n137), .Y(n312) );
  OR2X4 U1259 ( .A(n509), .B(n516), .Y(n983) );
  NAND2X2 U1260 ( .A(n379), .B(n388), .Y(n191) );
  INVX2 U1261 ( .A(n288), .Y(n286) );
  NAND2X1 U1262 ( .A(n334), .B(n297), .Y(n80) );
  NAND2X1 U1263 ( .A(n984), .B(n283), .Y(n77) );
  NAND2XL U1264 ( .A(n378), .B(n371), .Y(n184) );
  INVX2 U1265 ( .A(n105), .Y(n103) );
  INVX2 U1266 ( .A(n116), .Y(n114) );
  NAND2X1 U1267 ( .A(n988), .B(n989), .Y(n100) );
  NOR2X1 U1268 ( .A(n100), .B(n91), .Y(n89) );
  ADDFHX1 U1269 ( .A(n535), .B(n538), .CI(n533), .CO(n530), .S(n531) );
  NOR2X1 U1270 ( .A(n545), .B(n546), .Y(n296) );
  NAND2X1 U1271 ( .A(n342), .B(n341), .Y(n116) );
  NAND2XL U1272 ( .A(n346), .B(n343), .Y(n129) );
  OR2X1 U1273 ( .A(n342), .B(n341), .Y(n988) );
  OR2X1 U1274 ( .A(n340), .B(n339), .Y(n989) );
  INVX2 U1275 ( .A(n338), .Y(n339) );
  NAND2X1 U1276 ( .A(n340), .B(n339), .Y(n105) );
  NOR2X1 U1277 ( .A(n564), .B(n338), .Y(n91) );
  NAND2X1 U1278 ( .A(n564), .B(n338), .Y(n92) );
  OAI2BB1X1 U1279 ( .A0N(n22), .A1N(n24), .B0(n552), .Y(n628) );
  ADDFX1 U1280 ( .A(n569), .B(n368), .CI(n612), .CO(n360), .S(n361) );
  OAI2BB1X1 U1281 ( .A0N(n28), .A1N(n30), .B0(n551), .Y(n612) );
  INVX2 U1282 ( .A(n743), .Y(n551) );
  CLKINVXL U1283 ( .A(n386), .Y(n387) );
  OAI2BB1X1 U1284 ( .A0N(n9), .A1N(n12), .B0(n554), .Y(n660) );
  ADDFHX1 U1285 ( .A(n574), .B(n588), .CI(n616), .CO(n404), .S(n405) );
  ADDFHX1 U1286 ( .A(n645), .B(n589), .CI(n631), .CO(n418), .S(n419) );
  ADDFHX1 U1287 ( .A(n595), .B(n680), .CI(n609), .CO(n496), .S(n497) );
  ADDFHX1 U1288 ( .A(n639), .B(n958), .CI(n667), .CO(n512), .S(n513) );
  ADDFHX1 U1289 ( .A(n579), .B(n678), .CI(n593), .CO(n474), .S(n475) );
  ADDFHX1 U1290 ( .A(n627), .B(n684), .CI(n641), .CO(n528), .S(n529) );
  ADDFHX1 U1291 ( .A(n647), .B(n577), .CI(n605), .CO(n444), .S(n445) );
  OAI2BB1X1 U1292 ( .A0N(n867), .A1N(n6), .B0(n555), .Y(n676) );
  ADDFHX1 U1293 ( .A(n632), .B(n576), .CI(n618), .CO(n430), .S(n431) );
  ADDHXL U1294 ( .A(n679), .B(n650), .CO(n486), .S(n487) );
  OAI2BB1X1 U1295 ( .A0N(n34), .A1N(n36), .B0(n550), .Y(n596) );
  INVX2 U1296 ( .A(n726), .Y(n550) );
  ADDFX2 U1297 ( .A(n669), .B(n655), .CI(n534), .CO(n526), .S(n527) );
  ADDFX2 U1298 ( .A(n671), .B(n542), .CI(n539), .CO(n536), .S(n537) );
  ADDFX2 U1299 ( .A(n659), .B(n688), .CI(n673), .CO(n544), .S(n545) );
  NAND2BX1 U1300 ( .AN(b[0]), .B(n991), .Y(n827) );
  ADDFX2 U1301 ( .A(n566), .B(n345), .CI(n348), .CO(n342), .S(n343) );
  INVX2 U1302 ( .A(n344), .Y(n345) );
  CLKINVXL U1303 ( .A(n354), .Y(n355) );
  ADDFX2 U1304 ( .A(n344), .B(n565), .CI(n580), .CO(n340), .S(n341) );
  INVX2 U1305 ( .A(n709), .Y(n549) );
  INVX2 U1306 ( .A(n811), .Y(n555) );
  OAI2BB1X1 U1307 ( .A0N(n46), .A1N(n48), .B0(n548), .Y(n564) );
  INVX2 U1308 ( .A(n692), .Y(n548) );
  XOR2X1 U1309 ( .A(n995), .B(a[8]), .Y(n847) );
  BUFX12 U1310 ( .A(a[7]), .Y(n994) );
  XOR2X1 U1311 ( .A(n993), .B(a[4]), .Y(n849) );
  XOR2X1 U1312 ( .A(n992), .B(a[2]), .Y(n850) );
  BUFX12 U1313 ( .A(a[1]), .Y(n991) );
  XNOR2XL U1314 ( .A(b[15]), .B(n994), .Y(n760) );
  XNOR2XL U1315 ( .A(b[11]), .B(n991), .Y(n815) );
  XNOR2XL U1316 ( .A(b[14]), .B(n994), .Y(n761) );
  XNOR2XL U1317 ( .A(b[10]), .B(n991), .Y(n816) );
  XNOR2XL U1318 ( .A(b[14]), .B(n995), .Y(n744) );
  XNOR2XL U1319 ( .A(b[7]), .B(n991), .Y(n819) );
  XNOR2XL U1320 ( .A(b[14]), .B(n993), .Y(n778) );
  XNOR2XL U1321 ( .A(b[6]), .B(n991), .Y(n820) );
  XNOR2XL U1322 ( .A(b[11]), .B(n997), .Y(n713) );
  XNOR2XL U1323 ( .A(b[13]), .B(n995), .Y(n745) );
  XNOR2XL U1324 ( .A(b[6]), .B(n995), .Y(n752) );
  XNOR2XL U1325 ( .A(b[12]), .B(n996), .Y(n729) );
  XNOR2XL U1326 ( .A(b[10]), .B(n994), .Y(n765) );
  XNOR2XL U1327 ( .A(b[12]), .B(n995), .Y(n746) );
  XNOR2XL U1328 ( .A(b[5]), .B(n993), .Y(n787) );
  XNOR2XL U1329 ( .A(b[5]), .B(n995), .Y(n753) );
  XNOR2XL U1330 ( .A(b[15]), .B(n996), .Y(n726) );
  XNOR2XL U1331 ( .A(b[11]), .B(n996), .Y(n730) );
  XNOR2XL U1332 ( .A(b[10]), .B(n992), .Y(n799) );
  XNOR2XL U1333 ( .A(b[4]), .B(n991), .Y(n822) );
  XNOR2XL U1334 ( .A(b[7]), .B(n996), .Y(n734) );
  XNOR2XL U1335 ( .A(b[1]), .B(n996), .Y(n740) );
  XNOR2XL U1336 ( .A(b[12]), .B(n997), .Y(n712) );
  XNOR2XL U1337 ( .A(b[5]), .B(n996), .Y(n736) );
  XNOR2XL U1338 ( .A(b[11]), .B(n994), .Y(n764) );
  XNOR2XL U1339 ( .A(b[3]), .B(n991), .Y(n823) );
  XNOR2XL U1340 ( .A(b[6]), .B(n996), .Y(n735) );
  XNOR2XL U1341 ( .A(b[4]), .B(n996), .Y(n737) );
  XNOR2XL U1342 ( .A(b[8]), .B(n996), .Y(n733) );
  XNOR2XL U1343 ( .A(b[4]), .B(n993), .Y(n788) );
  XNOR2XL U1344 ( .A(b[10]), .B(n993), .Y(n782) );
  XNOR2XL U1345 ( .A(b[5]), .B(n991), .Y(n821) );
  XNOR2XL U1346 ( .A(b[8]), .B(n995), .Y(n750) );
  XNOR2XL U1347 ( .A(b[3]), .B(n993), .Y(n789) );
  XNOR2XL U1348 ( .A(b[1]), .B(n991), .Y(n825) );
  XNOR2XL U1349 ( .A(b[14]), .B(n996), .Y(n727) );
  XNOR2XL U1350 ( .A(b[6]), .B(n994), .Y(n769) );
  XNOR2XL U1351 ( .A(b[4]), .B(n994), .Y(n771) );
  XNOR2XL U1352 ( .A(b[3]), .B(n996), .Y(n738) );
  XNOR2XL U1353 ( .A(b[1]), .B(n995), .Y(n757) );
  XNOR2XL U1354 ( .A(b[7]), .B(n995), .Y(n751) );
  XNOR2XL U1355 ( .A(b[2]), .B(n993), .Y(n790) );
  XNOR2XL U1356 ( .A(b[2]), .B(n991), .Y(n824) );
  XNOR2XL U1357 ( .A(b[5]), .B(n994), .Y(n770) );
  XNOR2XL U1358 ( .A(b[3]), .B(n994), .Y(n772) );
  XNOR2XL U1359 ( .A(b[3]), .B(n995), .Y(n755) );
  XNOR2XL U1360 ( .A(b[4]), .B(n995), .Y(n754) );
  XNOR2XL U1361 ( .A(b[1]), .B(n993), .Y(n791) );
  XNOR2XL U1362 ( .A(b[6]), .B(n992), .Y(n803) );
  XNOR2XL U1363 ( .A(b[2]), .B(n994), .Y(n773) );
  XNOR2XL U1364 ( .A(b[7]), .B(n992), .Y(n802) );
  XNOR2XL U1365 ( .A(b[5]), .B(n992), .Y(n804) );
  XNOR2XL U1366 ( .A(b[13]), .B(n997), .Y(n711) );
  XNOR2XL U1367 ( .A(b[3]), .B(n992), .Y(n806) );
  XNOR2XL U1368 ( .A(b[4]), .B(n992), .Y(n805) );
  XNOR2XL U1369 ( .A(b[10]), .B(n995), .Y(n748) );
  XNOR2XL U1370 ( .A(b[10]), .B(n996), .Y(n731) );
  XNOR2XL U1371 ( .A(b[15]), .B(n997), .Y(n709) );
  XNOR2XL U1372 ( .A(b[2]), .B(n992), .Y(n807) );
  XNOR2XL U1373 ( .A(b[13]), .B(n996), .Y(n728) );
  XNOR2XL U1374 ( .A(b[8]), .B(n992), .Y(n801) );
  XNOR2XL U1375 ( .A(b[9]), .B(n995), .Y(n749) );
  XNOR2XL U1376 ( .A(b[11]), .B(n995), .Y(n747) );
  XNOR2XL U1377 ( .A(b[1]), .B(n992), .Y(n808) );
  XNOR2XL U1378 ( .A(b[14]), .B(n997), .Y(n710) );
  XNOR2XL U1379 ( .A(b[13]), .B(n998), .Y(n694) );
  XNOR2XL U1380 ( .A(b[14]), .B(n998), .Y(n693) );
  XNOR2XL U1381 ( .A(b[15]), .B(n998), .Y(n692) );
  OAI21XL U1382 ( .A0(n224), .A1(n216), .B0(n219), .Y(n215) );
  NOR2X4 U1383 ( .A(n211), .B(n216), .Y(n209) );
  OAI2BB1X1 U1384 ( .A0N(n40), .A1N(n42), .B0(n549), .Y(n580) );
  OAI22XL U1385 ( .A0(n42), .A1(n711), .B0(n710), .B1(n40), .Y(n581) );
  OAI22XL U1386 ( .A0(n42), .A1(n710), .B0(n709), .B1(n40), .Y(n344) );
  OAI22XL U1387 ( .A0(n42), .A1(n712), .B0(n711), .B1(n40), .Y(n582) );
  OAI22XL U1388 ( .A0(n42), .A1(n713), .B0(n712), .B1(n40), .Y(n583) );
  OAI22XL U1389 ( .A0(n42), .A1(n714), .B0(n713), .B1(n40), .Y(n584) );
  OAI22XL U1390 ( .A0(n42), .A1(n720), .B0(n719), .B1(n40), .Y(n590) );
  OAI22XL U1391 ( .A0(n42), .A1(n715), .B0(n714), .B1(n40), .Y(n585) );
  OAI22XL U1392 ( .A0(n42), .A1(n722), .B0(n721), .B1(n40), .Y(n592) );
  OAI22XL U1393 ( .A0(n42), .A1(n716), .B0(n715), .B1(n40), .Y(n586) );
  OAI22XL U1394 ( .A0(n42), .A1(n717), .B0(n716), .B1(n40), .Y(n587) );
  OAI22XL U1395 ( .A0(n42), .A1(n718), .B0(n717), .B1(n40), .Y(n588) );
  OAI22XL U1396 ( .A0(n42), .A1(n719), .B0(n718), .B1(n40), .Y(n589) );
  OAI22XL U1397 ( .A0(n42), .A1(n723), .B0(n722), .B1(n40), .Y(n593) );
  ADDHX1 U1398 ( .A(n683), .B(n654), .CO(n522), .S(n523) );
  OAI22XL U1399 ( .A0(n6), .A1(n818), .B0(n817), .B1(n867), .Y(n683) );
  NAND2BX1 U1400 ( .AN(b[0]), .B(n993), .Y(n793) );
  NOR2X4 U1401 ( .A(n241), .B(n238), .Y(n236) );
  INVX2 U1402 ( .A(n238), .Y(n324) );
  NAND2X1 U1403 ( .A(n690), .B(n675), .Y(n305) );
  NOR2X1 U1404 ( .A(n690), .B(n675), .Y(n304) );
  OAI2BB1X1 U1405 ( .A0N(n16), .A1N(n18), .B0(n553), .Y(n644) );
  OAI22XL U1406 ( .A0(n18), .A1(n785), .B0(n784), .B1(n16), .Y(n651) );
  OAI22XL U1407 ( .A0(n18), .A1(n783), .B0(n782), .B1(n16), .Y(n649) );
  OAI22XL U1408 ( .A0(n18), .A1(n791), .B0(n790), .B1(n16), .Y(n657) );
  OAI22XL U1409 ( .A0(n18), .A1(n779), .B0(n778), .B1(n16), .Y(n645) );
  OAI22XL U1410 ( .A0(n18), .A1(n787), .B0(n786), .B1(n16), .Y(n653) );
  OAI22XL U1411 ( .A0(n18), .A1(n781), .B0(n780), .B1(n16), .Y(n647) );
  OAI22XL U1412 ( .A0(n18), .A1(n789), .B0(n788), .B1(n16), .Y(n655) );
  ADDFHX1 U1413 ( .A(n560), .B(n642), .CI(n670), .CO(n532), .S(n533) );
  OAI21X2 U1414 ( .A0(n268), .A1(n256), .B0(n257), .Y(n255) );
  NOR2X4 U1415 ( .A(n423), .B(n436), .Y(n216) );
  ADDFX2 U1416 ( .A(n571), .B(n386), .CI(n628), .CO(n376), .S(n377) );
  NAND2BX1 U1417 ( .AN(b[0]), .B(n997), .Y(n725) );
  XNOR2X1 U1418 ( .A(b[0]), .B(n998), .Y(n707) );
  NOR2BXL U1419 ( .AN(b[0]), .B(n46), .Y(n579) );
  NOR2BXL U1420 ( .AN(b[0]), .B(n34), .Y(n611) );
  NOR2BXL U1421 ( .AN(b[0]), .B(n867), .Y(product[0]) );
  NOR2BXL U1422 ( .AN(b[0]), .B(n40), .Y(n595) );
  NOR2BXL U1423 ( .AN(b[0]), .B(n28), .Y(n627) );
  XNOR2X1 U1424 ( .A(b[0]), .B(n997), .Y(n724) );
  XNOR2X1 U1425 ( .A(b[0]), .B(n996), .Y(n741) );
  NOR2BXL U1426 ( .AN(b[0]), .B(n16), .Y(n659) );
  NAND2BX1 U1427 ( .AN(b[0]), .B(n995), .Y(n759) );
  XNOR2X1 U1428 ( .A(b[0]), .B(n995), .Y(n758) );
  NOR2BXL U1429 ( .AN(b[0]), .B(n9), .Y(n675) );
  XNOR2X1 U1430 ( .A(b[0]), .B(n993), .Y(n792) );
  XNOR2X1 U1431 ( .A(b[0]), .B(n992), .Y(n809) );
endmodule


module PE_DW_mult_tc_16 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n6, n9, n12, n16, n18, n22, n24, n30, n34, n36, n40, n42, n46, n48,
         n51, n52, n53, n55, n56, n57, n58, n59, n60, n62, n63, n64, n66, n67,
         n68, n69, n70, n72, n73, n75, n76, n77, n80, n81, n82, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n103, n105, n106, n107, n108, n109, n110, n114, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n140, n141,
         n142, n143, n144, n145, n148, n149, n151, n154, n155, n156, n157,
         n158, n159, n160, n164, n166, n167, n168, n169, n170, n171, n176,
         n177, n178, n181, n182, n183, n184, n185, n186, n187, n188, n191,
         n192, n193, n194, n196, n199, n200, n201, n203, n204, n205, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n219, n220,
         n221, n222, n224, n227, n228, n229, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n244, n245, n246, n247,
         n248, n249, n251, n254, n255, n256, n257, n259, n260, n261, n262,
         n264, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n281, n283, n284, n286, n288, n289, n290,
         n292, n294, n295, n296, n297, n298, n300, n302, n303, n304, n305,
         n307, n308, n311, n312, n313, n315, n318, n319, n320, n321, n323,
         n324, n325, n326, n327, n329, n330, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n844, n845, n846, n848, n849, n850, n851, n867, n868, n869, n870,
         n871, n872, n874, n875, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002;

  AOI21X1 U60 ( .A0(n123), .A1(n89), .B0(n90), .Y(n88) );
  AOI21X1 U72 ( .A0(n123), .A1(n98), .B0(n99), .Y(n97) );
  AOI21X1 U76 ( .A0(n114), .A1(n987), .B0(n103), .Y(n101) );
  AOI21X1 U106 ( .A0(n126), .A1(n151), .B0(n127), .Y(n125) );
  AOI21X1 U114 ( .A0(n953), .A1(n131), .B0(n132), .Y(n130) );
  AOI21X1 U118 ( .A0(n160), .A1(n135), .B0(n136), .Y(n134) );
  AOI21X1 U132 ( .A0(n160), .A1(n313), .B0(n151), .Y(n145) );
  AOI21X1 U144 ( .A0(n953), .A1(n155), .B0(n156), .Y(n154) );
  NOR2X2 U169 ( .A(n370), .B(n363), .Y(n170) );
  NOR2X2 U181 ( .A(n378), .B(n371), .Y(n183) );
  NOR2X2 U203 ( .A(n389), .B(n398), .Y(n199) );
  NOR2X2 U211 ( .A(n399), .B(n410), .Y(n204) );
  NOR2X2 U231 ( .A(n423), .B(n436), .Y(n216) );
  NOR2X2 U291 ( .A(n499), .B(n508), .Y(n260) );
  ADDFHX4 U389 ( .A(n392), .B(n390), .CI(n381), .CO(n378), .S(n379) );
  ADDFHX4 U394 ( .A(n402), .B(n400), .CI(n391), .CO(n388), .S(n389) );
  ADDFHX4 U399 ( .A(n403), .B(n412), .CI(n401), .CO(n398), .S(n399) );
  ADDFHX4 U411 ( .A(n427), .B(n438), .CI(n425), .CO(n422), .S(n423) );
  ADDFHX4 U414 ( .A(n590), .B(n448), .CI(n446), .CO(n428), .S(n429) );
  ADDFHX4 U418 ( .A(n441), .B(n452), .CI(n439), .CO(n436), .S(n437) );
  ADDFHX4 U445 ( .A(n493), .B(n500), .CI(n491), .CO(n488), .S(n489) );
  ADDFHX4 U455 ( .A(n513), .B(n518), .CI(n511), .CO(n508), .S(n509) );
  OAI22X1 U478 ( .A0(n48), .A1(n693), .B0(n692), .B1(n46), .Y(n338) );
  OAI22X1 U479 ( .A0(n48), .A1(n694), .B0(n693), .B1(n46), .Y(n565) );
  OAI22X1 U480 ( .A0(n48), .A1(n695), .B0(n694), .B1(n46), .Y(n566) );
  OAI22X1 U481 ( .A0(n48), .A1(n696), .B0(n695), .B1(n46), .Y(n567) );
  OAI22X1 U483 ( .A0(n48), .A1(n698), .B0(n697), .B1(n46), .Y(n569) );
  OAI22X1 U484 ( .A0(n48), .A1(n699), .B0(n698), .B1(n46), .Y(n570) );
  OAI22X1 U486 ( .A0(n48), .A1(n701), .B0(n700), .B1(n46), .Y(n572) );
  OAI22X1 U487 ( .A0(n48), .A1(n702), .B0(n701), .B1(n46), .Y(n573) );
  OAI22X1 U488 ( .A0(n48), .A1(n703), .B0(n702), .B1(n46), .Y(n574) );
  OAI22X1 U514 ( .A0(n42), .A1(n710), .B0(n709), .B1(n951), .Y(n344) );
  OAI22X1 U515 ( .A0(n42), .A1(n711), .B0(n710), .B1(n951), .Y(n581) );
  OAI22X1 U516 ( .A0(n42), .A1(n712), .B0(n711), .B1(n951), .Y(n582) );
  OAI22X1 U517 ( .A0(n42), .A1(n713), .B0(n712), .B1(n951), .Y(n583) );
  OAI22X1 U518 ( .A0(n42), .A1(n714), .B0(n713), .B1(n951), .Y(n584) );
  OAI22X1 U519 ( .A0(n42), .A1(n715), .B0(n714), .B1(n951), .Y(n585) );
  OAI22X1 U526 ( .A0(n42), .A1(n722), .B0(n721), .B1(n951), .Y(n592) );
  OAI22X1 U527 ( .A0(n42), .A1(n723), .B0(n722), .B1(n951), .Y(n593) );
  OAI22X1 U550 ( .A0(n36), .A1(n727), .B0(n726), .B1(n34), .Y(n354) );
  OAI22X1 U551 ( .A0(n36), .A1(n728), .B0(n727), .B1(n34), .Y(n597) );
  OAI22X1 U552 ( .A0(n36), .A1(n729), .B0(n728), .B1(n34), .Y(n598) );
  OAI22X1 U554 ( .A0(n36), .A1(n731), .B0(n730), .B1(n34), .Y(n600) );
  OAI22X1 U555 ( .A0(n36), .A1(n732), .B0(n731), .B1(n34), .Y(n601) );
  OAI22X1 U556 ( .A0(n36), .A1(n733), .B0(n732), .B1(n34), .Y(n602) );
  OAI22X1 U557 ( .A0(n36), .A1(n734), .B0(n733), .B1(n34), .Y(n603) );
  OAI22X1 U558 ( .A0(n36), .A1(n735), .B0(n734), .B1(n34), .Y(n604) );
  OAI22X1 U559 ( .A0(n36), .A1(n736), .B0(n735), .B1(n34), .Y(n605) );
  OAI22X1 U563 ( .A0(n36), .A1(n740), .B0(n739), .B1(n34), .Y(n609) );
  OAI22X1 U586 ( .A0(n30), .A1(n744), .B0(n743), .B1(n989), .Y(n368) );
  OAI22X1 U587 ( .A0(n30), .A1(n745), .B0(n744), .B1(n989), .Y(n613) );
  OAI22X1 U588 ( .A0(n30), .A1(n746), .B0(n745), .B1(n989), .Y(n614) );
  OAI22X1 U589 ( .A0(n30), .A1(n747), .B0(n746), .B1(n989), .Y(n615) );
  OAI22X1 U590 ( .A0(n30), .A1(n748), .B0(n747), .B1(n989), .Y(n616) );
  OAI22X1 U591 ( .A0(n30), .A1(n749), .B0(n748), .B1(n989), .Y(n617) );
  OAI22X1 U592 ( .A0(n30), .A1(n750), .B0(n749), .B1(n989), .Y(n618) );
  OAI22X1 U593 ( .A0(n30), .A1(n751), .B0(n750), .B1(n989), .Y(n619) );
  OAI22X1 U594 ( .A0(n30), .A1(n752), .B0(n751), .B1(n989), .Y(n620) );
  OAI22X1 U597 ( .A0(n30), .A1(n755), .B0(n754), .B1(n989), .Y(n623) );
  OAI22X1 U619 ( .A0(n24), .A1(n872), .B0(n22), .B1(n776), .Y(n560) );
  OAI22X1 U655 ( .A0(n18), .A1(n960), .B0(n956), .B1(n793), .Y(n561) );
  OAI22X1 U659 ( .A0(n18), .A1(n779), .B0(n778), .B1(n956), .Y(n645) );
  OAI22X1 U661 ( .A0(n18), .A1(n781), .B0(n780), .B1(n956), .Y(n647) );
  OAI22X1 U663 ( .A0(n18), .A1(n783), .B0(n782), .B1(n956), .Y(n649) );
  OAI22X1 U665 ( .A0(n18), .A1(n785), .B0(n784), .B1(n956), .Y(n651) );
  OAI22X1 U667 ( .A0(n18), .A1(n787), .B0(n786), .B1(n956), .Y(n653) );
  OAI22X1 U668 ( .A0(n18), .A1(n788), .B0(n787), .B1(n956), .Y(n654) );
  OAI22X1 U671 ( .A0(n18), .A1(n791), .B0(n790), .B1(n956), .Y(n657) );
  OAI22X1 U672 ( .A0(n18), .A1(n792), .B0(n791), .B1(n956), .Y(n658) );
  OAI22X1 U694 ( .A0(n12), .A1(n795), .B0(n794), .B1(n9), .Y(n434) );
  OAI22X1 U695 ( .A0(n12), .A1(n796), .B0(n795), .B1(n9), .Y(n661) );
  OAI22X1 U730 ( .A0(n6), .A1(n812), .B0(n811), .B1(n867), .Y(n677) );
  OAI22X1 U731 ( .A0(n6), .A1(n813), .B0(n812), .B1(n867), .Y(n678) );
  OAI22X1 U732 ( .A0(n6), .A1(n814), .B0(n813), .B1(n867), .Y(n679) );
  OAI22X1 U733 ( .A0(n6), .A1(n815), .B0(n814), .B1(n867), .Y(n680) );
  OAI22X1 U734 ( .A0(n6), .A1(n816), .B0(n815), .B1(n867), .Y(n681) );
  OAI22X1 U735 ( .A0(n6), .A1(n817), .B0(n816), .B1(n867), .Y(n682) );
  OAI22X1 U736 ( .A0(n6), .A1(n818), .B0(n817), .B1(n867), .Y(n683) );
  OAI22X1 U737 ( .A0(n6), .A1(n819), .B0(n818), .B1(n867), .Y(n684) );
  OAI22X1 U738 ( .A0(n6), .A1(n820), .B0(n819), .B1(n867), .Y(n685) );
  OAI22X1 U740 ( .A0(n6), .A1(n822), .B0(n821), .B1(n867), .Y(n687) );
  OAI22X1 U741 ( .A0(n6), .A1(n823), .B0(n822), .B1(n867), .Y(n688) );
  OAI22X1 U742 ( .A0(n6), .A1(n824), .B0(n823), .B1(n867), .Y(n689) );
  OAI22X1 U743 ( .A0(n6), .A1(n825), .B0(n824), .B1(n867), .Y(n690) );
  XNOR2X4 U788 ( .A(n999), .B(a[14]), .Y(n46) );
  XNOR2X4 U791 ( .A(n998), .B(a[12]), .Y(n40) );
  NAND2X4 U792 ( .A(n34), .B(n846), .Y(n36) );
  XNOR2X4 U794 ( .A(n997), .B(a[10]), .Y(n34) );
  NAND2X4 U798 ( .A(n22), .B(n848), .Y(n24) );
  NAND2X4 U801 ( .A(n955), .B(n849), .Y(n18) );
  XNOR2X4 U803 ( .A(n994), .B(a[4]), .Y(n16) );
  NAND2X4 U804 ( .A(n9), .B(n850), .Y(n12) );
  XNOR2X4 U806 ( .A(n993), .B(a[2]), .Y(n9) );
  NAND2X4 U807 ( .A(n851), .B(n867), .Y(n6) );
  ADDFHX2 U812 ( .A(n442), .B(n429), .CI(n440), .CO(n424), .S(n425) );
  AOI21X1 U813 ( .A0(n953), .A1(n193), .B0(n194), .Y(n192) );
  OAI22X1 U814 ( .A0(n24), .A1(n766), .B0(n765), .B1(n22), .Y(n633) );
  OR2X4 U815 ( .A(n547), .B(n674), .Y(n985) );
  ADDHX1 U816 ( .A(n683), .B(n654), .CO(n522), .S(n523) );
  ADDFHX1 U817 ( .A(n469), .B(n478), .CI(n467), .CO(n464), .S(n465) );
  CMPR32X1 U818 ( .A(n485), .B(n483), .C(n492), .CO(n478), .S(n479) );
  INVX3 U819 ( .A(n235), .Y(n234) );
  XOR2X4 U820 ( .A(n996), .B(a[8]), .Y(n988) );
  OAI21X2 U821 ( .A0(n242), .A1(n238), .B0(n239), .Y(n237) );
  XNOR2X2 U822 ( .A(n273), .B(n75), .Y(product[9]) );
  OAI22X2 U823 ( .A0(n30), .A1(n757), .B0(n756), .B1(n989), .Y(n625) );
  NAND2X2 U824 ( .A(n327), .B(n981), .Y(n256) );
  ADDFHX1 U825 ( .A(n559), .B(n626), .CI(n640), .CO(n520), .S(n521) );
  NAND2XL U826 ( .A(n953), .B(n186), .Y(n943) );
  INVX1 U827 ( .A(n187), .Y(n944) );
  AND2X4 U828 ( .A(n943), .B(n944), .Y(n185) );
  XOR2X4 U829 ( .A(n185), .B(n62), .Y(product[22]) );
  XOR3X4 U830 ( .A(n466), .B(n455), .C(n453), .Y(n451) );
  NAND2XL U831 ( .A(n453), .B(n466), .Y(n945) );
  NAND2X1 U832 ( .A(n455), .B(n466), .Y(n946) );
  NAND2XL U833 ( .A(n455), .B(n453), .Y(n947) );
  NAND3X1 U834 ( .A(n946), .B(n947), .C(n945), .Y(n450) );
  ADDFHX1 U835 ( .A(n472), .B(n470), .CI(n459), .CO(n454), .S(n455) );
  ADDFHX2 U836 ( .A(n482), .B(n471), .CI(n480), .CO(n466), .S(n467) );
  ADDFHX4 U837 ( .A(n461), .B(n457), .CI(n468), .CO(n452), .S(n453) );
  NAND2X1 U838 ( .A(n437), .B(n450), .Y(n228) );
  OR2X4 U839 ( .A(n30), .B(n754), .Y(n948) );
  OR2X4 U840 ( .A(n753), .B(n989), .Y(n949) );
  NAND2X4 U841 ( .A(n948), .B(n949), .Y(n622) );
  XNOR2XL U842 ( .A(b[4]), .B(n997), .Y(n754) );
  ADDFHX2 U843 ( .A(n622), .B(n958), .CI(n608), .CO(n482), .S(n483) );
  OAI22X2 U844 ( .A0(n6), .A1(n821), .B0(n820), .B1(n867), .Y(n686) );
  ADDFHX2 U845 ( .A(n557), .B(n664), .CI(n636), .CO(n484), .S(n485) );
  OAI22X2 U846 ( .A0(n42), .A1(n869), .B0(n951), .B1(n725), .Y(n557) );
  NOR2X2 U847 ( .A(n966), .B(n259), .Y(n257) );
  ADDFHX1 U848 ( .A(n637), .B(n665), .CI(n623), .CO(n494), .S(n495) );
  XNOR2XL U849 ( .A(b[2]), .B(n999), .Y(n722) );
  XNOR2XL U850 ( .A(b[2]), .B(n993), .Y(n824) );
  BUFX3 U851 ( .A(n40), .Y(n950) );
  BUFX8 U852 ( .A(n40), .Y(n951) );
  NOR2X2 U853 ( .A(n411), .B(n422), .Y(n211) );
  INVX4 U854 ( .A(n51), .Y(n952) );
  INVX8 U855 ( .A(n952), .Y(n953) );
  OAI21X2 U856 ( .A0(n207), .A1(n235), .B0(n208), .Y(n51) );
  AOI21X2 U857 ( .A0(n325), .A1(n251), .B0(n244), .Y(n242) );
  AOI21X2 U858 ( .A0(n209), .A1(n222), .B0(n210), .Y(n208) );
  ADDFHX1 U859 ( .A(n621), .B(n663), .CI(n649), .CO(n472), .S(n473) );
  INVX3 U860 ( .A(n16), .Y(n954) );
  CLKINVX2 U861 ( .A(n954), .Y(n955) );
  INVX12 U862 ( .A(n954), .Y(n956) );
  OAI22X1 U863 ( .A0(n42), .A1(n724), .B0(n723), .B1(n951), .Y(n594) );
  OAI22XL U864 ( .A0(n30), .A1(n756), .B0(n755), .B1(n989), .Y(n624) );
  OAI22XL U865 ( .A0(n30), .A1(n871), .B0(n989), .B1(n759), .Y(n559) );
  INVX3 U866 ( .A(n988), .Y(n989) );
  ADDFHX1 U867 ( .A(n558), .B(n610), .CI(n666), .CO(n504), .S(n505) );
  NAND2XL U868 ( .A(n325), .B(n326), .Y(n241) );
  NOR2X2 U869 ( .A(n465), .B(n476), .Y(n238) );
  XNOR2X2 U870 ( .A(n953), .B(n970), .Y(product[19]) );
  OAI22X2 U871 ( .A0(n18), .A1(n786), .B0(n785), .B1(n956), .Y(n652) );
  ADDFHX1 U872 ( .A(n635), .B(n607), .CI(n486), .CO(n470), .S(n471) );
  OAI22XL U873 ( .A0(n36), .A1(n738), .B0(n737), .B1(n34), .Y(n607) );
  ADDFHX1 U874 ( .A(n604), .B(n646), .CI(n435), .CO(n432), .S(n433) );
  OAI22X2 U875 ( .A0(n42), .A1(n721), .B0(n720), .B1(n951), .Y(n591) );
  XNOR2X2 U876 ( .A(b[14]), .B(n994), .Y(n795) );
  XNOR2X2 U877 ( .A(b[14]), .B(n993), .Y(n812) );
  XNOR2X2 U878 ( .A(b[15]), .B(n994), .Y(n794) );
  XNOR2X2 U879 ( .A(b[15]), .B(n993), .Y(n811) );
  INVX1 U880 ( .A(n594), .Y(n957) );
  CLKINVX2 U881 ( .A(n957), .Y(n958) );
  XNOR2X1 U882 ( .A(b[3]), .B(n999), .Y(n721) );
  XNOR2X1 U883 ( .A(b[3]), .B(n997), .Y(n755) );
  XNOR2X1 U884 ( .A(b[3]), .B(n996), .Y(n772) );
  XNOR2X1 U885 ( .A(b[3]), .B(n1000), .Y(n704) );
  ADDFHX1 U886 ( .A(n595), .B(n680), .CI(n609), .CO(n496), .S(n497) );
  XNOR2X2 U887 ( .A(b[8]), .B(n996), .Y(n767) );
  XNOR2X1 U888 ( .A(b[8]), .B(n995), .Y(n784) );
  XNOR2XL U889 ( .A(b[8]), .B(n993), .Y(n818) );
  XNOR2X2 U890 ( .A(b[8]), .B(n997), .Y(n750) );
  XNOR2X1 U891 ( .A(b[8]), .B(n994), .Y(n801) );
  XNOR2X1 U892 ( .A(b[7]), .B(n995), .Y(n785) );
  XNOR2X1 U893 ( .A(b[7]), .B(n998), .Y(n734) );
  XNOR2X2 U894 ( .A(b[7]), .B(n996), .Y(n768) );
  XNOR2X1 U895 ( .A(b[7]), .B(n997), .Y(n751) );
  XNOR2XL U896 ( .A(b[7]), .B(n993), .Y(n819) );
  XNOR2X2 U897 ( .A(b[9]), .B(n996), .Y(n766) );
  XNOR2X1 U898 ( .A(b[9]), .B(n995), .Y(n783) );
  XNOR2XL U899 ( .A(b[9]), .B(n993), .Y(n817) );
  XNOR2X2 U900 ( .A(b[9]), .B(n994), .Y(n800) );
  OAI22X2 U901 ( .A0(n48), .A1(n706), .B0(n705), .B1(n46), .Y(n577) );
  OAI22XL U902 ( .A0(n48), .A1(n700), .B0(n699), .B1(n46), .Y(n571) );
  NAND2X4 U903 ( .A(n46), .B(n844), .Y(n48) );
  XNOR2X2 U904 ( .A(b[10]), .B(n996), .Y(n765) );
  XNOR2X2 U905 ( .A(b[10]), .B(n994), .Y(n799) );
  XNOR2X2 U906 ( .A(b[10]), .B(n993), .Y(n816) );
  XNOR2X1 U907 ( .A(b[10]), .B(n995), .Y(n782) );
  XNOR2X1 U908 ( .A(b[13]), .B(n995), .Y(n779) );
  XNOR2XL U909 ( .A(b[13]), .B(n993), .Y(n813) );
  XNOR2X2 U910 ( .A(b[13]), .B(n994), .Y(n796) );
  XNOR2X1 U911 ( .A(b[4]), .B(n998), .Y(n737) );
  XNOR2X2 U912 ( .A(b[4]), .B(n996), .Y(n771) );
  XNOR2X1 U913 ( .A(b[4]), .B(n995), .Y(n788) );
  XNOR2X2 U914 ( .A(b[4]), .B(n1000), .Y(n703) );
  NAND2X4 U915 ( .A(n950), .B(n845), .Y(n42) );
  XNOR2X2 U916 ( .A(b[11]), .B(n993), .Y(n815) );
  XNOR2X2 U917 ( .A(b[11]), .B(n994), .Y(n798) );
  XNOR2X1 U918 ( .A(b[11]), .B(n995), .Y(n781) );
  XNOR2X1 U919 ( .A(b[11]), .B(n996), .Y(n764) );
  BUFX8 U920 ( .A(a[11]), .Y(n998) );
  BUFX8 U921 ( .A(a[13]), .Y(n999) );
  INVX2 U922 ( .A(n245), .Y(n325) );
  NOR2X1 U923 ( .A(n477), .B(n488), .Y(n245) );
  CMPR32X1 U924 ( .A(n584), .B(n570), .C(n369), .CO(n366), .S(n367) );
  ADDFX2 U925 ( .A(n582), .B(n568), .CI(n355), .CO(n352), .S(n353) );
  ADDFX2 U926 ( .A(n354), .B(n567), .CI(n596), .CO(n348), .S(n349) );
  NAND2X2 U927 ( .A(n451), .B(n464), .Y(n233) );
  NOR2X2 U928 ( .A(n437), .B(n450), .Y(n227) );
  NAND2X1 U929 ( .A(n411), .B(n422), .Y(n212) );
  ADDFHX1 U930 ( .A(n382), .B(n373), .CI(n380), .CO(n370), .S(n371) );
  NOR2X1 U931 ( .A(n241), .B(n238), .Y(n236) );
  OR2XL U932 ( .A(n24), .B(n775), .Y(n968) );
  NAND2X1 U933 ( .A(n964), .B(n965), .Y(n562) );
  ADDHXL U934 ( .A(n681), .B(n652), .CO(n506), .S(n507) );
  ADDHXL U935 ( .A(n679), .B(n650), .CO(n486), .S(n487) );
  INVX2 U936 ( .A(n266), .Y(n264) );
  ADDFX1 U937 ( .A(n647), .B(n577), .CI(n605), .CO(n444), .S(n445) );
  CMPR32X1 U938 ( .A(n585), .B(n599), .C(n613), .CO(n374), .S(n375) );
  ADDFX1 U939 ( .A(n586), .B(n614), .CI(n387), .CO(n384), .S(n385) );
  AOI21X1 U940 ( .A0(n269), .A1(n277), .B0(n270), .Y(n268) );
  ADDFX2 U941 ( .A(n597), .B(n583), .CI(n366), .CO(n358), .S(n359) );
  ADDFX2 U942 ( .A(n361), .B(n359), .CI(n364), .CO(n356), .S(n357) );
  NOR2X1 U943 ( .A(n356), .B(n351), .Y(n148) );
  ADDFHX1 U944 ( .A(n415), .B(n424), .CI(n413), .CO(n410), .S(n411) );
  NAND2XL U945 ( .A(n324), .B(n239), .Y(n70) );
  NAND2X2 U946 ( .A(n399), .B(n410), .Y(n205) );
  INVX2 U947 ( .A(n166), .Y(n164) );
  ADDFX2 U948 ( .A(n360), .B(n353), .CI(n358), .CO(n350), .S(n351) );
  NAND2X1 U949 ( .A(n356), .B(n351), .Y(n149) );
  ADDFX2 U950 ( .A(n581), .B(n352), .CI(n349), .CO(n346), .S(n347) );
  NAND2XL U951 ( .A(n122), .B(n98), .Y(n96) );
  NOR2X1 U952 ( .A(n204), .B(n199), .Y(n193) );
  NOR2BXL U953 ( .AN(n193), .B(n188), .Y(n186) );
  NAND2X1 U954 ( .A(n370), .B(n363), .Y(n171) );
  INVX2 U955 ( .A(n53), .Y(n177) );
  NOR2X1 U956 ( .A(n350), .B(n347), .Y(n137) );
  NOR2X1 U957 ( .A(n53), .B(n144), .Y(n142) );
  NOR2X1 U958 ( .A(n346), .B(n343), .Y(n128) );
  NOR2X1 U959 ( .A(n53), .B(n96), .Y(n94) );
  NAND2X2 U960 ( .A(n193), .B(n181), .Y(n53) );
  NAND2X1 U961 ( .A(n209), .B(n221), .Y(n207) );
  NOR2X2 U962 ( .A(n211), .B(n216), .Y(n209) );
  OR2X1 U963 ( .A(n12), .B(n874), .Y(n964) );
  NAND2X1 U964 ( .A(n968), .B(n969), .Y(n642) );
  ADDFX2 U965 ( .A(n639), .B(n653), .CI(n667), .CO(n512), .S(n513) );
  ADDFX2 U966 ( .A(n668), .B(n523), .CI(n528), .CO(n518), .S(n519) );
  ADDFX2 U967 ( .A(n522), .B(n515), .CI(n520), .CO(n510), .S(n511) );
  ADDFX2 U968 ( .A(n638), .B(n624), .CI(n507), .CO(n502), .S(n503) );
  ADDFHX1 U969 ( .A(n514), .B(n512), .CI(n505), .CO(n500), .S(n501) );
  XOR2X2 U970 ( .A(n993), .B(a[0]), .Y(n851) );
  ADDFX2 U971 ( .A(n651), .B(n506), .CI(n497), .CO(n492), .S(n493) );
  NAND2X1 U972 ( .A(n509), .B(n516), .Y(n266) );
  ADDFHX1 U973 ( .A(n504), .B(n502), .CI(n495), .CO(n490), .S(n491) );
  ADDFX2 U974 ( .A(n487), .B(n496), .CI(n494), .CO(n480), .S(n481) );
  ADDFX2 U975 ( .A(n662), .B(n606), .CI(n620), .CO(n458), .S(n459) );
  ADDFX2 U976 ( .A(n634), .B(n463), .CI(n474), .CO(n456), .S(n457) );
  ADDFX2 U977 ( .A(n462), .B(n449), .CI(n460), .CO(n442), .S(n443) );
  XNOR2X1 U978 ( .A(n990), .B(n591), .Y(n449) );
  ADDFX2 U979 ( .A(n475), .B(n484), .CI(n473), .CO(n468), .S(n469) );
  NOR2X1 U980 ( .A(n489), .B(n498), .Y(n248) );
  ADDFX2 U981 ( .A(n617), .B(n603), .CI(n432), .CO(n416), .S(n417) );
  ADDFHX1 U982 ( .A(n481), .B(n490), .CI(n479), .CO(n476), .S(n477) );
  ADDFHX1 U983 ( .A(n428), .B(n417), .CI(n426), .CO(n412), .S(n413) );
  ADDFX2 U984 ( .A(n430), .B(n421), .CI(n419), .CO(n414), .S(n415) );
  ADDFHX1 U985 ( .A(n444), .B(n433), .CI(n431), .CO(n426), .S(n427) );
  ADDFHX1 U986 ( .A(n458), .B(n447), .CI(n445), .CO(n440), .S(n441) );
  ADDFHX1 U987 ( .A(n456), .B(n443), .CI(n454), .CO(n438), .S(n439) );
  ADDFX2 U988 ( .A(n418), .B(n416), .CI(n414), .CO(n400), .S(n401) );
  ADDFX2 U989 ( .A(n420), .B(n405), .CI(n407), .CO(n402), .S(n403) );
  ADDFX2 U990 ( .A(n615), .B(n406), .CI(n404), .CO(n392), .S(n393) );
  ADDFX2 U991 ( .A(n395), .B(n397), .CI(n393), .CO(n390), .S(n391) );
  ADDFX2 U992 ( .A(n598), .B(n376), .CI(n374), .CO(n364), .S(n365) );
  ADDFX2 U993 ( .A(n384), .B(n377), .CI(n375), .CO(n372), .S(n373) );
  ADDFX2 U994 ( .A(n394), .B(n385), .CI(n383), .CO(n380), .S(n381) );
  NOR2X1 U995 ( .A(n137), .B(n128), .Y(n126) );
  OAI21X2 U996 ( .A0(n268), .A1(n256), .B0(n257), .Y(n255) );
  INVX2 U997 ( .A(n261), .Y(n259) );
  NAND2X1 U998 ( .A(n465), .B(n476), .Y(n239) );
  INVX2 U999 ( .A(a[0]), .Y(n867) );
  NAND2X1 U1000 ( .A(n321), .B(n219), .Y(n67) );
  ADDFX2 U1001 ( .A(n367), .B(n365), .CI(n372), .CO(n362), .S(n363) );
  NOR2X1 U1002 ( .A(n53), .B(n170), .Y(n168) );
  NOR2X1 U1003 ( .A(n227), .B(n232), .Y(n221) );
  OAI21X1 U1004 ( .A0(n211), .A1(n219), .B0(n212), .Y(n210) );
  OAI21X2 U1005 ( .A0(n227), .A1(n233), .B0(n228), .Y(n222) );
  NOR2X1 U1006 ( .A(n53), .B(n120), .Y(n118) );
  NOR2X1 U1007 ( .A(n53), .B(n109), .Y(n107) );
  XOR2X1 U1008 ( .A(n213), .B(n66), .Y(product[18]) );
  NAND2X1 U1009 ( .A(n320), .B(n212), .Y(n66) );
  NOR2X1 U1010 ( .A(n967), .B(n215), .Y(n213) );
  XOR2X1 U1011 ( .A(n201), .B(n64), .Y(product[20]) );
  XOR2X1 U1012 ( .A(n192), .B(n63), .Y(product[21]) );
  XOR2X1 U1013 ( .A(n154), .B(n59), .Y(product[25]) );
  XNOR2X1 U1014 ( .A(n176), .B(n978), .Y(product[23]) );
  XOR2X1 U1015 ( .A(n141), .B(n58), .Y(product[26]) );
  XOR2X1 U1016 ( .A(n130), .B(n57), .Y(product[27]) );
  INVX2 U1017 ( .A(n91), .Y(n308) );
  NOR2X1 U1018 ( .A(n53), .B(n87), .Y(n85) );
  AND2X1 U1019 ( .A(n975), .B(n307), .Y(product[1]) );
  BUFX8 U1020 ( .A(a[5]), .Y(n995) );
  XOR2X1 U1021 ( .A(n229), .B(n68), .Y(product[16]) );
  AOI21X1 U1022 ( .A0(n234), .A1(n323), .B0(n231), .Y(n229) );
  OAI22X1 U1023 ( .A0(n12), .A1(n799), .B0(n798), .B1(n9), .Y(n664) );
  ADDHX1 U1024 ( .A(n689), .B(n562), .CO(n546), .S(n547) );
  XOR2X1 U1025 ( .A(n220), .B(n67), .Y(product[17]) );
  ADDFHX2 U1026 ( .A(n503), .B(n510), .CI(n501), .CO(n498), .S(n499) );
  AND2X2 U1027 ( .A(n214), .B(n234), .Y(n967) );
  ADDFX2 U1028 ( .A(n682), .B(n611), .CI(n625), .CO(n514), .S(n515) );
  AOI21X1 U1029 ( .A0(n234), .A1(n221), .B0(n222), .Y(n220) );
  INVX3 U1030 ( .A(n255), .Y(n254) );
  INVX2 U1031 ( .A(n260), .Y(n327) );
  NAND2X1 U1032 ( .A(n995), .B(a[6]), .Y(n962) );
  NAND2X4 U1033 ( .A(n960), .B(n961), .Y(n963) );
  NAND2X4 U1034 ( .A(n962), .B(n963), .Y(n22) );
  INVX2 U1035 ( .A(n995), .Y(n960) );
  INVX1 U1036 ( .A(a[6]), .Y(n961) );
  OAI22XL U1037 ( .A0(n24), .A1(n774), .B0(n773), .B1(n22), .Y(n641) );
  OAI22XL U1038 ( .A0(n24), .A1(n771), .B0(n770), .B1(n22), .Y(n638) );
  OAI22XL U1039 ( .A0(n24), .A1(n768), .B0(n767), .B1(n22), .Y(n635) );
  OAI22XL U1040 ( .A0(n24), .A1(n767), .B0(n766), .B1(n22), .Y(n634) );
  OAI22XL U1041 ( .A0(n24), .A1(n764), .B0(n763), .B1(n22), .Y(n631) );
  OAI22XL U1042 ( .A0(n24), .A1(n772), .B0(n771), .B1(n22), .Y(n639) );
  OAI22XL U1043 ( .A0(n24), .A1(n773), .B0(n772), .B1(n22), .Y(n640) );
  OAI22XL U1044 ( .A0(n24), .A1(n765), .B0(n764), .B1(n22), .Y(n632) );
  OAI22XL U1045 ( .A0(n24), .A1(n769), .B0(n768), .B1(n22), .Y(n636) );
  OAI22XL U1046 ( .A0(n24), .A1(n763), .B0(n762), .B1(n22), .Y(n630) );
  OAI22XL U1047 ( .A0(n24), .A1(n761), .B0(n760), .B1(n22), .Y(n386) );
  OAI22XL U1048 ( .A0(n24), .A1(n762), .B0(n761), .B1(n22), .Y(n629) );
  OR2X1 U1049 ( .A(n9), .B(n810), .Y(n965) );
  AND2X4 U1050 ( .A(n327), .B(n264), .Y(n966) );
  INVX4 U1051 ( .A(n1002), .Y(n1001) );
  XNOR2XL U1052 ( .A(b[1]), .B(n996), .Y(n774) );
  OR2X1 U1053 ( .A(n774), .B(n22), .Y(n969) );
  XNOR2XL U1054 ( .A(n1001), .B(n996), .Y(n775) );
  OAI21X2 U1055 ( .A0(n183), .A1(n191), .B0(n184), .Y(n182) );
  XOR2X1 U1056 ( .A(n996), .B(a[6]), .Y(n848) );
  NAND2X2 U1057 ( .A(n159), .B(n313), .Y(n144) );
  NAND2X1 U1058 ( .A(n315), .B(n980), .Y(n157) );
  NAND2XL U1059 ( .A(n159), .B(n135), .Y(n133) );
  CMPR32X1 U1060 ( .A(n535), .B(n538), .C(n533), .CO(n530), .S(n531) );
  ADDFX1 U1061 ( .A(n521), .B(n526), .CI(n519), .CO(n516), .S(n517) );
  NAND2X1 U1062 ( .A(n319), .B(n205), .Y(n970) );
  CLKINVXL U1063 ( .A(n232), .Y(n323) );
  INVX2 U1064 ( .A(n248), .Y(n326) );
  NAND2BX1 U1065 ( .AN(n188), .B(n191), .Y(n63) );
  NAND2XL U1066 ( .A(n980), .B(n166), .Y(n60) );
  NAND2X1 U1067 ( .A(n389), .B(n398), .Y(n200) );
  INVX2 U1068 ( .A(n148), .Y(n313) );
  NAND2X1 U1069 ( .A(n499), .B(n508), .Y(n261) );
  INVX1 U1070 ( .A(n283), .Y(n281) );
  NAND2BX1 U1071 ( .AN(n304), .B(n305), .Y(n82) );
  NAND2X1 U1072 ( .A(n362), .B(n357), .Y(n166) );
  NAND2XL U1073 ( .A(n122), .B(n986), .Y(n109) );
  ADDFHX1 U1074 ( .A(n560), .B(n642), .CI(n670), .CO(n532), .S(n533) );
  OAI22XL U1075 ( .A0(n30), .A1(n758), .B0(n757), .B1(n989), .Y(n626) );
  ADDHX1 U1076 ( .A(n677), .B(n648), .CO(n462), .S(n463) );
  CLKINVXL U1077 ( .A(n794), .Y(n554) );
  ADDFX2 U1078 ( .A(n574), .B(n588), .CI(n616), .CO(n404), .S(n405) );
  ADDFHX1 U1079 ( .A(n573), .B(n408), .CI(n644), .CO(n396), .S(n397) );
  XOR2X1 U1080 ( .A(n999), .B(a[12]), .Y(n845) );
  XNOR2XL U1081 ( .A(b[6]), .B(n997), .Y(n752) );
  XNOR2XL U1082 ( .A(b[6]), .B(n996), .Y(n769) );
  XNOR2XL U1083 ( .A(b[5]), .B(n997), .Y(n753) );
  XNOR2XL U1084 ( .A(b[5]), .B(n998), .Y(n736) );
  XNOR2XL U1085 ( .A(b[6]), .B(n998), .Y(n735) );
  XNOR2XL U1086 ( .A(b[6]), .B(n999), .Y(n718) );
  XNOR2XL U1087 ( .A(b[5]), .B(n999), .Y(n719) );
  XNOR2XL U1088 ( .A(b[8]), .B(n1000), .Y(n699) );
  XNOR2XL U1089 ( .A(b[7]), .B(n1000), .Y(n700) );
  XNOR2XL U1090 ( .A(b[12]), .B(n1000), .Y(n695) );
  XNOR2X1 U1091 ( .A(n240), .B(n70), .Y(product[14]) );
  NAND2BX1 U1092 ( .AN(n227), .B(n228), .Y(n68) );
  OAI21XL U1093 ( .A0(n992), .A1(n144), .B0(n145), .Y(n143) );
  XOR2X1 U1094 ( .A(n262), .B(n73), .Y(product[11]) );
  XOR2X1 U1095 ( .A(n247), .B(n971), .Y(product[13]) );
  AND2X1 U1096 ( .A(n325), .B(n246), .Y(n971) );
  CLKINVXL U1097 ( .A(n277), .Y(n276) );
  NAND2XL U1098 ( .A(n329), .B(n272), .Y(n75) );
  OAI21XL U1099 ( .A0(n276), .A1(n274), .B0(n275), .Y(n273) );
  CLKINVXL U1100 ( .A(n271), .Y(n329) );
  NAND2BX1 U1101 ( .AN(n183), .B(n184), .Y(n62) );
  XOR2X1 U1102 ( .A(n276), .B(n76), .Y(product[8]) );
  NAND2XL U1103 ( .A(n330), .B(n275), .Y(n76) );
  CLKINVXL U1104 ( .A(n274), .Y(n330) );
  XOR2X1 U1105 ( .A(n167), .B(n60), .Y(product[24]) );
  BUFX8 U1106 ( .A(n52), .Y(n992) );
  CLKINVXL U1107 ( .A(n290), .Y(n289) );
  CLKINVX4 U1108 ( .A(n980), .Y(n977) );
  NAND2X1 U1109 ( .A(n313), .B(n126), .Y(n124) );
  INVX2 U1110 ( .A(n149), .Y(n151) );
  NAND2XL U1111 ( .A(n122), .B(n89), .Y(n87) );
  NAND2XL U1112 ( .A(n982), .B(n983), .Y(n278) );
  INVX1 U1113 ( .A(n288), .Y(n286) );
  NAND2XL U1114 ( .A(n477), .B(n488), .Y(n246) );
  NAND2XL U1115 ( .A(n982), .B(n283), .Y(n77) );
  AOI21XL U1116 ( .A0(n289), .A1(n983), .B0(n286), .Y(n284) );
  NAND2XL U1117 ( .A(n312), .B(n140), .Y(n58) );
  XOR2X1 U1118 ( .A(n972), .B(n289), .Y(product[6]) );
  AND2X1 U1119 ( .A(n983), .B(n288), .Y(n972) );
  NAND2XL U1120 ( .A(n985), .B(n302), .Y(n81) );
  NAND2BX1 U1121 ( .AN(n296), .B(n297), .Y(n80) );
  XOR2X1 U1122 ( .A(n106), .B(n55), .Y(product[29]) );
  XOR2XL U1123 ( .A(n973), .B(n295), .Y(product[5]) );
  AND2X1 U1124 ( .A(n984), .B(n294), .Y(n973) );
  XOR2X1 U1125 ( .A(n117), .B(n56), .Y(product[28]) );
  OAI21XL U1126 ( .A0(n158), .A1(n124), .B0(n125), .Y(n123) );
  AOI21X1 U1127 ( .A0(n123), .A1(n986), .B0(n114), .Y(n110) );
  XOR2X1 U1128 ( .A(n93), .B(n974), .Y(product[30]) );
  NAND2X1 U1129 ( .A(n308), .B(n92), .Y(n974) );
  NAND2XL U1130 ( .A(n531), .B(n536), .Y(n283) );
  ADDFX1 U1131 ( .A(n529), .B(n532), .CI(n527), .CO(n524), .S(n525) );
  NAND2XL U1132 ( .A(n547), .B(n674), .Y(n302) );
  OR2XL U1133 ( .A(n691), .B(n563), .Y(n975) );
  ADDFHX1 U1134 ( .A(n643), .B(n686), .CI(n657), .CO(n538), .S(n539) );
  ADDFX1 U1135 ( .A(n671), .B(n542), .CI(n539), .CO(n536), .S(n537) );
  OAI22XL U1136 ( .A0(n18), .A1(n790), .B0(n789), .B1(n956), .Y(n656) );
  OAI22XL U1137 ( .A0(n18), .A1(n789), .B0(n788), .B1(n956), .Y(n655) );
  ADDFX1 U1138 ( .A(n561), .B(n672), .CI(n543), .CO(n540), .S(n541) );
  CLKINVXL U1139 ( .A(n994), .Y(n874) );
  XNOR2XL U1140 ( .A(n1001), .B(n995), .Y(n792) );
  ADDFX1 U1141 ( .A(n659), .B(n688), .CI(n673), .CO(n544), .S(n545) );
  CMPR32X1 U1142 ( .A(n579), .B(n678), .C(n593), .CO(n474), .S(n475) );
  OAI22XL U1143 ( .A0(n36), .A1(n739), .B0(n738), .B1(n34), .Y(n608) );
  OAI22XL U1144 ( .A0(n24), .A1(n770), .B0(n769), .B1(n22), .Y(n637) );
  OAI22XL U1145 ( .A0(n42), .A1(n720), .B0(n719), .B1(n951), .Y(n590) );
  XNOR2XL U1146 ( .A(n1001), .B(n994), .Y(n809) );
  OAI22XL U1147 ( .A0(n48), .A1(n707), .B0(n706), .B1(n46), .Y(n578) );
  ADDFHX1 U1148 ( .A(n602), .B(n630), .CI(n991), .CO(n406), .S(n407) );
  OAI22XL U1149 ( .A0(n48), .A1(n704), .B0(n703), .B1(n46), .Y(n575) );
  CLKINVXL U1150 ( .A(n993), .Y(n875) );
  NAND2BXL U1151 ( .AN(n1001), .B(n993), .Y(n827) );
  NAND2BXL U1152 ( .AN(b[0]), .B(n994), .Y(n810) );
  NAND2BX1 U1153 ( .AN(b[0]), .B(n999), .Y(n725) );
  OAI22XL U1154 ( .A0(n18), .A1(n782), .B0(n781), .B1(n956), .Y(n648) );
  OAI22XL U1155 ( .A0(n48), .A1(n705), .B0(n704), .B1(n46), .Y(n576) );
  NAND2BXL U1156 ( .AN(b[0]), .B(n995), .Y(n793) );
  OAI22XL U1157 ( .A0(n42), .A1(n719), .B0(n718), .B1(n951), .Y(n589) );
  OAI22XL U1158 ( .A0(n42), .A1(n718), .B0(n717), .B1(n951), .Y(n588) );
  CLKINVXL U1159 ( .A(n996), .Y(n872) );
  CLKINVXL U1160 ( .A(n777), .Y(n553) );
  CLKINVXL U1161 ( .A(n997), .Y(n871) );
  CLKINVXL U1162 ( .A(n999), .Y(n869) );
  CLKINVXL U1163 ( .A(n760), .Y(n552) );
  OAI22XL U1164 ( .A0(n42), .A1(n717), .B0(n716), .B1(n951), .Y(n587) );
  OAI22XL U1165 ( .A0(n42), .A1(n716), .B0(n715), .B1(n951), .Y(n586) );
  OAI22XL U1166 ( .A0(n36), .A1(n730), .B0(n729), .B1(n34), .Y(n599) );
  CLKINVXL U1167 ( .A(n743), .Y(n551) );
  ADDFX1 U1168 ( .A(n569), .B(n368), .CI(n612), .CO(n360), .S(n361) );
  OAI22XL U1169 ( .A0(n48), .A1(n697), .B0(n696), .B1(n46), .Y(n568) );
  XNOR2X1 U1170 ( .A(b[2]), .B(n997), .Y(n756) );
  NAND2BX4 U1171 ( .AN(n988), .B(n976), .Y(n30) );
  XOR2X2 U1172 ( .A(n997), .B(a[8]), .Y(n976) );
  XNOR2X1 U1173 ( .A(b[2]), .B(n994), .Y(n807) );
  XNOR2X1 U1174 ( .A(b[2]), .B(n996), .Y(n773) );
  XNOR2X1 U1175 ( .A(b[2]), .B(n998), .Y(n739) );
  XNOR2X1 U1176 ( .A(b[2]), .B(n1000), .Y(n705) );
  BUFX12 U1177 ( .A(a[15]), .Y(n1000) );
  XNOR2X1 U1178 ( .A(b[1]), .B(n1000), .Y(n706) );
  XNOR2X1 U1179 ( .A(b[5]), .B(n1000), .Y(n702) );
  XNOR2X1 U1180 ( .A(b[6]), .B(n1000), .Y(n701) );
  XNOR2XL U1181 ( .A(b[15]), .B(n1000), .Y(n692) );
  INVX2 U1182 ( .A(n122), .Y(n120) );
  NOR2X1 U1183 ( .A(n157), .B(n124), .Y(n122) );
  NAND2X1 U1184 ( .A(n318), .B(n200), .Y(n64) );
  CLKINVXL U1185 ( .A(n199), .Y(n318) );
  CLKINVXL U1186 ( .A(n216), .Y(n321) );
  CLKINVXL U1187 ( .A(n211), .Y(n320) );
  CLKINVXL U1188 ( .A(n238), .Y(n324) );
  XNOR2X2 U1189 ( .A(n234), .B(n69), .Y(product[15]) );
  NAND2XL U1190 ( .A(n323), .B(n233), .Y(n69) );
  INVX2 U1191 ( .A(n268), .Y(n267) );
  INVX2 U1192 ( .A(n992), .Y(n178) );
  CLKINVXL U1193 ( .A(n222), .Y(n224) );
  INVX2 U1194 ( .A(n158), .Y(n160) );
  NOR2XL U1195 ( .A(n53), .B(n133), .Y(n131) );
  INVX2 U1196 ( .A(n157), .Y(n159) );
  NOR2BXL U1197 ( .AN(n221), .B(n216), .Y(n214) );
  CLKINVXL U1198 ( .A(n204), .Y(n319) );
  CLKINVXL U1199 ( .A(n233), .Y(n231) );
  CLKINVXL U1200 ( .A(n205), .Y(n203) );
  OAI21XL U1201 ( .A0(n992), .A1(n96), .B0(n97), .Y(n95) );
  INVX2 U1202 ( .A(n101), .Y(n99) );
  AOI2BB1X4 U1203 ( .A0N(n977), .A1N(n171), .B0(n164), .Y(n158) );
  INVX2 U1204 ( .A(n170), .Y(n315) );
  OAI21XL U1205 ( .A0(n992), .A1(n87), .B0(n88), .Y(n86) );
  OAI21XL U1206 ( .A0(n992), .A1(n170), .B0(n171), .Y(n169) );
  NOR2X2 U1207 ( .A(n188), .B(n183), .Y(n181) );
  INVX2 U1208 ( .A(n249), .Y(n251) );
  INVX2 U1209 ( .A(n246), .Y(n244) );
  NAND2X1 U1210 ( .A(n313), .B(n149), .Y(n59) );
  NOR2XL U1211 ( .A(n53), .B(n157), .Y(n155) );
  OAI21X1 U1212 ( .A0(n271), .A1(n275), .B0(n272), .Y(n270) );
  NOR2X1 U1213 ( .A(n271), .B(n274), .Y(n269) );
  NOR2X2 U1214 ( .A(n451), .B(n464), .Y(n232) );
  NAND2XL U1215 ( .A(n327), .B(n261), .Y(n73) );
  AOI21X1 U1216 ( .A0(n267), .A1(n981), .B0(n264), .Y(n262) );
  AND2X1 U1217 ( .A(n315), .B(n171), .Y(n978) );
  OAI21X1 U1218 ( .A0(n254), .A1(n248), .B0(n249), .Y(n247) );
  OAI21XL U1219 ( .A0(n196), .A1(n188), .B0(n191), .Y(n187) );
  CLKINVXL U1220 ( .A(n194), .Y(n196) );
  NAND2X2 U1221 ( .A(n423), .B(n436), .Y(n219) );
  XOR2X1 U1222 ( .A(n254), .B(n72), .Y(product[12]) );
  NAND2XL U1223 ( .A(n326), .B(n249), .Y(n72) );
  OAI21XL U1224 ( .A0(n992), .A1(n120), .B0(n121), .Y(n119) );
  INVX2 U1225 ( .A(n123), .Y(n121) );
  XOR2X1 U1226 ( .A(n267), .B(n979), .Y(product[10]) );
  AND2X1 U1227 ( .A(n981), .B(n266), .Y(n979) );
  INVX2 U1228 ( .A(n100), .Y(n98) );
  OAI21XL U1229 ( .A0(n140), .A1(n128), .B0(n129), .Y(n127) );
  OR2X4 U1230 ( .A(n362), .B(n357), .Y(n980) );
  OAI21X1 U1231 ( .A0(n101), .A1(n91), .B0(n92), .Y(n90) );
  NOR2X1 U1232 ( .A(n517), .B(n524), .Y(n271) );
  OAI21X1 U1233 ( .A0(n278), .A1(n290), .B0(n279), .Y(n277) );
  AOI21X1 U1234 ( .A0(n982), .A1(n286), .B0(n281), .Y(n279) );
  NAND2X2 U1235 ( .A(n379), .B(n388), .Y(n191) );
  NOR2X1 U1236 ( .A(n525), .B(n530), .Y(n274) );
  CLKINVXL U1237 ( .A(n137), .Y(n312) );
  NAND2X1 U1238 ( .A(n987), .B(n105), .Y(n55) );
  OAI21XL U1239 ( .A0(n992), .A1(n109), .B0(n110), .Y(n108) );
  NAND2X2 U1240 ( .A(n489), .B(n498), .Y(n249) );
  NAND2X1 U1241 ( .A(n311), .B(n129), .Y(n57) );
  CLKINVXL U1242 ( .A(n128), .Y(n311) );
  OAI21XL U1243 ( .A0(n992), .A1(n133), .B0(n134), .Y(n132) );
  OAI21XL U1244 ( .A0(n149), .A1(n137), .B0(n140), .Y(n136) );
  NAND2X1 U1245 ( .A(n517), .B(n524), .Y(n272) );
  NAND2XL U1246 ( .A(n378), .B(n371), .Y(n184) );
  NAND2X1 U1247 ( .A(n525), .B(n530), .Y(n275) );
  OR2X4 U1248 ( .A(n509), .B(n516), .Y(n981) );
  NAND2X1 U1249 ( .A(n986), .B(n116), .Y(n56) );
  AOI21X1 U1250 ( .A0(n295), .A1(n984), .B0(n292), .Y(n290) );
  INVX2 U1251 ( .A(n294), .Y(n292) );
  XOR2X1 U1252 ( .A(n284), .B(n77), .Y(product[7]) );
  OAI21X1 U1253 ( .A0(n298), .A1(n296), .B0(n297), .Y(n295) );
  OAI21X1 U1254 ( .A0(n304), .A1(n307), .B0(n305), .Y(n303) );
  AOI21X1 U1255 ( .A0(n985), .A1(n303), .B0(n300), .Y(n298) );
  INVX2 U1256 ( .A(n302), .Y(n300) );
  INVX2 U1257 ( .A(n105), .Y(n103) );
  INVX2 U1258 ( .A(n116), .Y(n114) );
  NOR2X1 U1259 ( .A(n148), .B(n137), .Y(n135) );
  NAND2X1 U1260 ( .A(n986), .B(n987), .Y(n100) );
  NOR2X1 U1261 ( .A(n100), .B(n91), .Y(n89) );
  OR2X1 U1262 ( .A(n531), .B(n536), .Y(n982) );
  NAND2X1 U1263 ( .A(n350), .B(n347), .Y(n140) );
  OR2X1 U1264 ( .A(n537), .B(n540), .Y(n983) );
  OR2X1 U1265 ( .A(n541), .B(n544), .Y(n984) );
  NAND2X1 U1266 ( .A(n691), .B(n563), .Y(n307) );
  NAND2X1 U1267 ( .A(n537), .B(n540), .Y(n288) );
  NAND2XL U1268 ( .A(n346), .B(n343), .Y(n129) );
  NOR2X1 U1269 ( .A(n545), .B(n546), .Y(n296) );
  NOR2X1 U1270 ( .A(n690), .B(n675), .Y(n304) );
  NAND2X1 U1271 ( .A(n541), .B(n544), .Y(n294) );
  NAND2X1 U1272 ( .A(n342), .B(n341), .Y(n116) );
  NAND2XL U1273 ( .A(n690), .B(n675), .Y(n305) );
  NAND2X1 U1274 ( .A(n545), .B(n546), .Y(n297) );
  OR2X1 U1275 ( .A(n342), .B(n341), .Y(n986) );
  OR2X1 U1276 ( .A(n340), .B(n339), .Y(n987) );
  INVX2 U1277 ( .A(n338), .Y(n339) );
  NAND2X1 U1278 ( .A(n340), .B(n339), .Y(n105) );
  NOR2X1 U1279 ( .A(n564), .B(n338), .Y(n91) );
  NAND2X1 U1280 ( .A(n564), .B(n338), .Y(n92) );
  OAI2BB1X1 U1281 ( .A0N(n34), .A1N(n36), .B0(n550), .Y(n596) );
  INVX2 U1282 ( .A(n726), .Y(n550) );
  OAI2BB1X1 U1283 ( .A0N(n22), .A1N(n24), .B0(n552), .Y(n628) );
  CLKINVXL U1284 ( .A(n434), .Y(n435) );
  ADDFHX1 U1285 ( .A(n632), .B(n576), .CI(n618), .CO(n430), .S(n431) );
  NOR2BXL U1286 ( .AN(n1001), .B(n46), .Y(n579) );
  ADDFX2 U1287 ( .A(n566), .B(n345), .CI(n348), .CO(n342), .S(n343) );
  INVX1 U1288 ( .A(n344), .Y(n345) );
  OAI22XL U1289 ( .A0(n48), .A1(n868), .B0(n46), .B1(n708), .Y(n556) );
  BUFX2 U1290 ( .A(n633), .Y(n990) );
  OAI22XL U1291 ( .A0(n36), .A1(n741), .B0(n740), .B1(n34), .Y(n610) );
  OAI22XL U1292 ( .A0(n36), .A1(n870), .B0(n34), .B1(n742), .Y(n558) );
  INVX1 U1293 ( .A(n368), .Y(n369) );
  OAI22XL U1294 ( .A0(n30), .A1(n753), .B0(n752), .B1(n989), .Y(n621) );
  ADDFHX1 U1295 ( .A(n645), .B(n589), .CI(n631), .CO(n418), .S(n419) );
  OAI2BB1X1 U1296 ( .A0N(n956), .A1N(n18), .B0(n553), .Y(n644) );
  CMPR32X1 U1297 ( .A(n600), .B(n572), .C(n396), .CO(n382), .S(n383) );
  ADDFHX1 U1298 ( .A(n669), .B(n655), .CI(n534), .CO(n526), .S(n527) );
  ADDHXL U1299 ( .A(n685), .B(n656), .CO(n534), .S(n535) );
  NOR2BXL U1300 ( .AN(n1001), .B(n951), .Y(n595) );
  ADDFHX1 U1301 ( .A(n629), .B(n587), .CI(n601), .CO(n394), .S(n395) );
  CLKINVXL U1302 ( .A(n354), .Y(n355) );
  ADDFX2 U1303 ( .A(n619), .B(n661), .CI(n676), .CO(n446), .S(n447) );
  OAI2BB1X1 U1304 ( .A0N(n867), .A1N(n6), .B0(n555), .Y(n676) );
  CLKINVXL U1305 ( .A(n386), .Y(n387) );
  OAI2BB1X1 U1306 ( .A0N(n989), .A1N(n30), .B0(n551), .Y(n612) );
  OR2X1 U1307 ( .A(n990), .B(n591), .Y(n448) );
  ADDFHX1 U1308 ( .A(n627), .B(n684), .CI(n641), .CO(n528), .S(n529) );
  NOR2BXL U1309 ( .AN(n1001), .B(n989), .Y(n627) );
  NOR2BXL U1310 ( .AN(n1001), .B(n34), .Y(n611) );
  XNOR2X1 U1311 ( .A(n1001), .B(n1000), .Y(n707) );
  INVX2 U1312 ( .A(b[0]), .Y(n1002) );
  NOR2BXL U1313 ( .AN(n1001), .B(n22), .Y(n643) );
  NAND2BX1 U1314 ( .AN(b[0]), .B(n1000), .Y(n708) );
  ADDHXL U1315 ( .A(n687), .B(n658), .CO(n542), .S(n543) );
  NAND2BXL U1316 ( .AN(n1001), .B(n996), .Y(n776) );
  NAND2BX1 U1317 ( .AN(n1001), .B(n997), .Y(n759) );
  XNOR2X1 U1318 ( .A(n1001), .B(n999), .Y(n724) );
  NAND2BX1 U1319 ( .AN(n1001), .B(n998), .Y(n742) );
  XNOR2X1 U1320 ( .A(n1001), .B(n998), .Y(n741) );
  NOR2BXL U1321 ( .AN(n1001), .B(n956), .Y(n659) );
  OAI22XL U1322 ( .A0(n6), .A1(n826), .B0(n825), .B1(n867), .Y(n691) );
  ADDFX2 U1323 ( .A(n344), .B(n565), .CI(n580), .CO(n340), .S(n341) );
  OAI2BB1X1 U1324 ( .A0N(n951), .A1N(n42), .B0(n549), .Y(n580) );
  INVX2 U1325 ( .A(n709), .Y(n549) );
  CLKINVXL U1326 ( .A(n811), .Y(n555) );
  INVX2 U1327 ( .A(n1000), .Y(n868) );
  INVX2 U1328 ( .A(n998), .Y(n870) );
  NOR2BXL U1329 ( .AN(n1001), .B(n867), .Y(product[0]) );
  OAI2BB1X1 U1330 ( .A0N(n46), .A1N(n48), .B0(n548), .Y(n564) );
  INVX2 U1331 ( .A(n692), .Y(n548) );
  XOR2X1 U1332 ( .A(n998), .B(a[10]), .Y(n846) );
  BUFX12 U1333 ( .A(a[9]), .Y(n997) );
  XOR2X1 U1334 ( .A(a[14]), .B(n1000), .Y(n844) );
  XOR2X1 U1335 ( .A(n995), .B(a[4]), .Y(n849) );
  BUFX12 U1336 ( .A(a[3]), .Y(n994) );
  XOR2X1 U1337 ( .A(n994), .B(a[2]), .Y(n850) );
  BUFX16 U1338 ( .A(a[1]), .Y(n993) );
  BUFX12 U1339 ( .A(a[7]), .Y(n996) );
  XNOR2XL U1340 ( .A(b[12]), .B(n994), .Y(n797) );
  XNOR2XL U1341 ( .A(b[15]), .B(n998), .Y(n726) );
  XNOR2XL U1342 ( .A(b[15]), .B(n996), .Y(n760) );
  XNOR2XL U1343 ( .A(b[15]), .B(n997), .Y(n743) );
  XNOR2XL U1344 ( .A(b[14]), .B(n998), .Y(n727) );
  XNOR2XL U1345 ( .A(b[14]), .B(n997), .Y(n744) );
  XNOR2XL U1346 ( .A(b[14]), .B(n996), .Y(n761) );
  XNOR2XL U1347 ( .A(b[12]), .B(n995), .Y(n780) );
  XNOR2XL U1348 ( .A(b[5]), .B(n995), .Y(n787) );
  XNOR2XL U1349 ( .A(b[13]), .B(n996), .Y(n762) );
  XNOR2XL U1350 ( .A(b[6]), .B(n995), .Y(n786) );
  XNOR2XL U1351 ( .A(b[9]), .B(n998), .Y(n732) );
  XNOR2XL U1352 ( .A(b[15]), .B(n995), .Y(n777) );
  XNOR2XL U1353 ( .A(b[3]), .B(n995), .Y(n789) );
  XNOR2XL U1354 ( .A(b[12]), .B(n996), .Y(n763) );
  XNOR2XL U1355 ( .A(b[7]), .B(n999), .Y(n717) );
  XNOR2XL U1356 ( .A(b[8]), .B(n998), .Y(n733) );
  XNOR2XL U1357 ( .A(b[4]), .B(n999), .Y(n720) );
  XNOR2XL U1358 ( .A(b[5]), .B(n996), .Y(n770) );
  XNOR2XL U1359 ( .A(b[1]), .B(n999), .Y(n723) );
  XNOR2XL U1360 ( .A(b[2]), .B(n995), .Y(n790) );
  XNOR2XL U1361 ( .A(b[3]), .B(n998), .Y(n738) );
  XNOR2XL U1362 ( .A(b[6]), .B(n994), .Y(n803) );
  XNOR2XL U1363 ( .A(b[3]), .B(n994), .Y(n806) );
  XNOR2XL U1364 ( .A(b[14]), .B(n995), .Y(n778) );
  XNOR2XL U1365 ( .A(b[1]), .B(n998), .Y(n740) );
  XNOR2XL U1366 ( .A(b[8]), .B(n999), .Y(n716) );
  XNOR2X1 U1367 ( .A(b[11]), .B(n1000), .Y(n696) );
  XNOR2XL U1368 ( .A(b[5]), .B(n994), .Y(n804) );
  XNOR2X1 U1369 ( .A(b[9]), .B(n1000), .Y(n698) );
  XNOR2XL U1370 ( .A(b[1]), .B(n994), .Y(n808) );
  XNOR2XL U1371 ( .A(b[1]), .B(n997), .Y(n757) );
  XNOR2XL U1372 ( .A(b[7]), .B(n994), .Y(n802) );
  XNOR2XL U1373 ( .A(b[11]), .B(n999), .Y(n713) );
  XNOR2XL U1374 ( .A(b[13]), .B(n997), .Y(n745) );
  XNOR2X1 U1375 ( .A(b[10]), .B(n1000), .Y(n697) );
  XNOR2XL U1376 ( .A(b[9]), .B(n999), .Y(n715) );
  XNOR2XL U1377 ( .A(b[12]), .B(n998), .Y(n729) );
  XNOR2XL U1378 ( .A(b[10]), .B(n999), .Y(n714) );
  XNOR2XL U1379 ( .A(b[12]), .B(n997), .Y(n746) );
  XNOR2XL U1380 ( .A(b[4]), .B(n994), .Y(n805) );
  XNOR2XL U1381 ( .A(b[13]), .B(n999), .Y(n711) );
  XNOR2XL U1382 ( .A(b[11]), .B(n998), .Y(n730) );
  XNOR2XL U1383 ( .A(b[12]), .B(n999), .Y(n712) );
  XNOR2XL U1384 ( .A(b[1]), .B(n995), .Y(n791) );
  XNOR2XL U1385 ( .A(b[10]), .B(n997), .Y(n748) );
  XNOR2XL U1386 ( .A(b[9]), .B(n997), .Y(n749) );
  XNOR2XL U1387 ( .A(b[11]), .B(n997), .Y(n747) );
  XNOR2XL U1388 ( .A(b[10]), .B(n998), .Y(n731) );
  XNOR2XL U1389 ( .A(b[15]), .B(n999), .Y(n709) );
  XNOR2XL U1390 ( .A(b[14]), .B(n999), .Y(n710) );
  XNOR2XL U1391 ( .A(b[13]), .B(n998), .Y(n728) );
  XNOR2XL U1392 ( .A(b[13]), .B(n1000), .Y(n694) );
  XNOR2XL U1393 ( .A(b[14]), .B(n1000), .Y(n693) );
  OAI22XL U1394 ( .A0(n18), .A1(n780), .B0(n779), .B1(n956), .Y(n646) );
  OAI22XL U1395 ( .A0(n36), .A1(n737), .B0(n736), .B1(n34), .Y(n606) );
  INVX2 U1396 ( .A(n408), .Y(n991) );
  OAI22XL U1397 ( .A0(n18), .A1(n778), .B0(n777), .B1(n956), .Y(n408) );
  OAI22XL U1398 ( .A0(n18), .A1(n784), .B0(n783), .B1(n956), .Y(n650) );
  XNOR2X1 U1399 ( .A(b[4]), .B(n993), .Y(n822) );
  XNOR2X1 U1400 ( .A(n1001), .B(n993), .Y(n826) );
  XNOR2X1 U1401 ( .A(b[12]), .B(n993), .Y(n814) );
  XNOR2X1 U1402 ( .A(b[3]), .B(n993), .Y(n823) );
  XNOR2X1 U1403 ( .A(b[6]), .B(n993), .Y(n820) );
  XNOR2X1 U1404 ( .A(b[1]), .B(n993), .Y(n825) );
  XNOR2X1 U1405 ( .A(b[5]), .B(n993), .Y(n821) );
  NOR2BX1 U1406 ( .AN(n1001), .B(n9), .Y(n675) );
  OAI22X1 U1407 ( .A0(n6), .A1(n875), .B0(n827), .B1(n867), .Y(n563) );
  OAI21X2 U1408 ( .A0(n199), .A1(n205), .B0(n200), .Y(n194) );
  XNOR2X1 U1409 ( .A(n1001), .B(n997), .Y(n758) );
  OAI22X1 U1410 ( .A0(n12), .A1(n809), .B0(n808), .B1(n9), .Y(n674) );
  OAI21XL U1411 ( .A0(n254), .A1(n241), .B0(n242), .Y(n240) );
  ADDFHX1 U1412 ( .A(n556), .B(n578), .CI(n592), .CO(n460), .S(n461) );
  AOI21X4 U1413 ( .A0(n255), .A1(n236), .B0(n237), .Y(n235) );
  OAI21XL U1414 ( .A0(n224), .A1(n216), .B0(n219), .Y(n215) );
  OAI21XL U1415 ( .A0(n992), .A1(n157), .B0(n158), .Y(n156) );
  ADDFX2 U1416 ( .A(n571), .B(n386), .CI(n628), .CO(n376), .S(n377) );
  ADDFX2 U1417 ( .A(n575), .B(n434), .CI(n660), .CO(n420), .S(n421) );
  OAI22XL U1418 ( .A0(n12), .A1(n802), .B0(n801), .B1(n9), .Y(n667) );
  OAI22XL U1419 ( .A0(n12), .A1(n806), .B0(n805), .B1(n9), .Y(n671) );
  OAI2BB1X1 U1420 ( .A0N(n9), .A1N(n12), .B0(n554), .Y(n660) );
  OAI22XL U1421 ( .A0(n12), .A1(n801), .B0(n800), .B1(n9), .Y(n666) );
  OAI22XL U1422 ( .A0(n12), .A1(n803), .B0(n802), .B1(n9), .Y(n668) );
  OAI22XL U1423 ( .A0(n12), .A1(n804), .B0(n803), .B1(n9), .Y(n669) );
  OAI22XL U1424 ( .A0(n12), .A1(n805), .B0(n804), .B1(n9), .Y(n670) );
  OAI22XL U1425 ( .A0(n12), .A1(n808), .B0(n807), .B1(n9), .Y(n673) );
  OAI22XL U1426 ( .A0(n12), .A1(n800), .B0(n799), .B1(n9), .Y(n665) );
  OAI22XL U1427 ( .A0(n12), .A1(n807), .B0(n806), .B1(n9), .Y(n672) );
  OAI22XL U1428 ( .A0(n12), .A1(n798), .B0(n797), .B1(n9), .Y(n663) );
  OAI22XL U1429 ( .A0(n12), .A1(n797), .B0(n796), .B1(n9), .Y(n662) );
  AOI21X1 U1430 ( .A0(n953), .A1(n177), .B0(n178), .Y(n176) );
  NOR2X4 U1431 ( .A(n379), .B(n388), .Y(n188) );
  AOI21XL U1432 ( .A0(n953), .A1(n85), .B0(n86), .Y(product[31]) );
  AOI21XL U1433 ( .A0(n953), .A1(n94), .B0(n95), .Y(n93) );
  AOI21XL U1434 ( .A0(n953), .A1(n118), .B0(n119), .Y(n117) );
  AOI21XL U1435 ( .A0(n953), .A1(n107), .B0(n108), .Y(n106) );
  AOI21XL U1436 ( .A0(n953), .A1(n319), .B0(n203), .Y(n201) );
  AOI21XL U1437 ( .A0(n953), .A1(n168), .B0(n169), .Y(n167) );
  AOI21XL U1438 ( .A0(n953), .A1(n142), .B0(n143), .Y(n141) );
  XNOR2X1 U1439 ( .A(n81), .B(n303), .Y(product[3]) );
  XOR2X1 U1440 ( .A(n82), .B(n307), .Y(product[2]) );
  XOR2X1 U1441 ( .A(n80), .B(n298), .Y(product[4]) );
  AOI21X4 U1442 ( .A0(n194), .A1(n181), .B0(n182), .Y(n52) );
endmodule


module PE_DW_mult_tc_19 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n6, n9, n12, n16, n18, n22, n24, n28, n30, n34, n36, n40, n42, n46,
         n48, n51, n52, n53, n55, n56, n57, n61, n62, n63, n64, n66, n67, n68,
         n70, n72, n73, n75, n76, n77, n80, n81, n82, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n103,
         n105, n106, n107, n108, n109, n110, n114, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n140, n141, n142, n143,
         n144, n145, n148, n149, n151, n154, n155, n156, n157, n158, n159,
         n160, n164, n165, n166, n167, n168, n169, n170, n171, n176, n177,
         n181, n182, n183, n184, n185, n186, n187, n188, n191, n192, n193,
         n194, n196, n199, n200, n201, n203, n204, n205, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n219, n220, n221, n222,
         n224, n227, n228, n229, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n244, n246, n247, n248, n249, n251,
         n254, n255, n256, n257, n259, n260, n261, n262, n264, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n281, n283, n284, n286, n288, n289, n290, n292, n294, n295,
         n296, n297, n298, n300, n302, n303, n304, n305, n307, n308, n312,
         n313, n314, n315, n319, n320, n321, n322, n323, n324, n326, n327,
         n329, n330, n334, n336, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n844,
         n845, n846, n847, n848, n849, n850, n851, n867, n868, n869, n870,
         n871, n872, n873, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009;

  AOI21X1 U60 ( .A0(n123), .A1(n89), .B0(n90), .Y(n88) );
  AOI21X1 U72 ( .A0(n123), .A1(n98), .B0(n99), .Y(n97) );
  AOI21X1 U76 ( .A0(n114), .A1(n998), .B0(n103), .Y(n101) );
  AOI21X1 U88 ( .A0(n123), .A1(n999), .B0(n114), .Y(n110) );
  AOI21X1 U118 ( .A0(n160), .A1(n135), .B0(n136), .Y(n134) );
  AOI21X1 U132 ( .A0(n160), .A1(n313), .B0(n151), .Y(n145) );
  NAND2X4 U175 ( .A(n193), .B(n181), .Y(n53) );
  NOR2X2 U199 ( .A(n204), .B(n199), .Y(n193) );
  NOR2X2 U211 ( .A(n399), .B(n410), .Y(n204) );
  NOR2X2 U256 ( .A(n241), .B(n238), .Y(n236) );
  NAND2X4 U281 ( .A(n489), .B(n498), .Y(n249) );
  AOI21X1 U286 ( .A0(n327), .A1(n264), .B0(n259), .Y(n257) );
  ADDFHX4 U378 ( .A(n361), .B(n359), .CI(n364), .CO(n356), .S(n357) );
  ADDFHX4 U385 ( .A(n382), .B(n373), .CI(n380), .CO(n370), .S(n371) );
  ADDFHX4 U389 ( .A(n392), .B(n390), .CI(n381), .CO(n378), .S(n379) );
  ADDFHX4 U394 ( .A(n402), .B(n400), .CI(n391), .CO(n388), .S(n389) );
  ADDFHX4 U399 ( .A(n403), .B(n412), .CI(n401), .CO(n398), .S(n399) );
  ADDFHX4 U405 ( .A(n415), .B(n424), .CI(n413), .CO(n410), .S(n411) );
  ADDFHX4 U426 ( .A(n455), .B(n466), .CI(n453), .CO(n450), .S(n451) );
  ADDFHX4 U439 ( .A(n481), .B(n490), .CI(n479), .CO(n476), .S(n477) );
  ADDFHX4 U445 ( .A(n493), .B(n500), .CI(n491), .CO(n488), .S(n489) );
  ADDFHX4 U450 ( .A(n503), .B(n510), .CI(n501), .CO(n498), .S(n499) );
  OAI22X1 U475 ( .A0(n48), .A1(n868), .B0(n46), .B1(n708), .Y(n556) );
  OAI22X1 U478 ( .A0(n48), .A1(n693), .B0(n692), .B1(n46), .Y(n338) );
  OAI22X1 U479 ( .A0(n48), .A1(n694), .B0(n693), .B1(n46), .Y(n565) );
  OAI22X1 U480 ( .A0(n48), .A1(n695), .B0(n694), .B1(n46), .Y(n566) );
  OAI22X1 U481 ( .A0(n48), .A1(n696), .B0(n695), .B1(n46), .Y(n567) );
  OAI22X1 U483 ( .A0(n48), .A1(n698), .B0(n697), .B1(n46), .Y(n569) );
  OAI22X1 U484 ( .A0(n48), .A1(n699), .B0(n698), .B1(n46), .Y(n570) );
  OAI22X1 U485 ( .A0(n48), .A1(n700), .B0(n699), .B1(n46), .Y(n571) );
  OAI22X1 U487 ( .A0(n48), .A1(n702), .B0(n701), .B1(n46), .Y(n573) );
  OAI22X1 U488 ( .A0(n48), .A1(n703), .B0(n702), .B1(n46), .Y(n574) );
  OAI22X1 U489 ( .A0(n48), .A1(n704), .B0(n703), .B1(n46), .Y(n575) );
  OAI22X1 U490 ( .A0(n48), .A1(n705), .B0(n704), .B1(n46), .Y(n576) );
  OAI22X1 U491 ( .A0(n48), .A1(n706), .B0(n705), .B1(n46), .Y(n577) );
  OAI22X1 U514 ( .A0(n42), .A1(n710), .B0(n709), .B1(n961), .Y(n344) );
  OAI22X1 U515 ( .A0(n42), .A1(n711), .B0(n710), .B1(n962), .Y(n581) );
  OAI22X1 U516 ( .A0(n42), .A1(n712), .B0(n711), .B1(n961), .Y(n582) );
  OAI22X1 U517 ( .A0(n42), .A1(n713), .B0(n712), .B1(n962), .Y(n583) );
  OAI22X1 U519 ( .A0(n42), .A1(n715), .B0(n714), .B1(n962), .Y(n585) );
  OAI22X1 U522 ( .A0(n42), .A1(n718), .B0(n717), .B1(n961), .Y(n588) );
  OAI22X1 U525 ( .A0(n42), .A1(n721), .B0(n720), .B1(n962), .Y(n591) );
  OAI22X1 U526 ( .A0(n42), .A1(n722), .B0(n721), .B1(n962), .Y(n592) );
  OAI22X1 U527 ( .A0(n42), .A1(n723), .B0(n722), .B1(n962), .Y(n593) );
  OAI22X1 U586 ( .A0(n30), .A1(n744), .B0(n743), .B1(n958), .Y(n368) );
  OAI22X1 U587 ( .A0(n30), .A1(n745), .B0(n744), .B1(n958), .Y(n613) );
  OAI22X1 U588 ( .A0(n30), .A1(n746), .B0(n745), .B1(n958), .Y(n614) );
  OAI22X1 U589 ( .A0(n30), .A1(n747), .B0(n746), .B1(n958), .Y(n615) );
  OAI22X1 U590 ( .A0(n30), .A1(n748), .B0(n747), .B1(n958), .Y(n616) );
  OAI22X1 U591 ( .A0(n30), .A1(n749), .B0(n748), .B1(n958), .Y(n617) );
  OAI22X1 U592 ( .A0(n30), .A1(n750), .B0(n749), .B1(n958), .Y(n618) );
  OAI22X1 U593 ( .A0(n30), .A1(n751), .B0(n750), .B1(n958), .Y(n619) );
  OAI22X1 U594 ( .A0(n30), .A1(n752), .B0(n751), .B1(n958), .Y(n620) );
  OAI22X1 U596 ( .A0(n30), .A1(n754), .B0(n753), .B1(n958), .Y(n622) );
  OAI22X1 U597 ( .A0(n30), .A1(n755), .B0(n754), .B1(n958), .Y(n623) );
  OAI22X1 U599 ( .A0(n30), .A1(n757), .B0(n756), .B1(n958), .Y(n625) );
  OAI22X1 U600 ( .A0(n30), .A1(n758), .B0(n757), .B1(n958), .Y(n626) );
  OAI22X1 U623 ( .A0(n24), .A1(n762), .B0(n761), .B1(n22), .Y(n629) );
  OAI22X1 U625 ( .A0(n24), .A1(n764), .B0(n763), .B1(n22), .Y(n631) );
  OAI22X1 U627 ( .A0(n24), .A1(n766), .B0(n765), .B1(n22), .Y(n633) );
  OAI22X1 U628 ( .A0(n24), .A1(n767), .B0(n766), .B1(n22), .Y(n634) );
  OAI22X1 U630 ( .A0(n24), .A1(n769), .B0(n768), .B1(n22), .Y(n636) );
  OAI22X1 U631 ( .A0(n24), .A1(n770), .B0(n769), .B1(n22), .Y(n637) );
  OAI22X1 U632 ( .A0(n24), .A1(n771), .B0(n770), .B1(n22), .Y(n638) );
  OAI22X1 U633 ( .A0(n24), .A1(n772), .B0(n771), .B1(n22), .Y(n639) );
  OAI22X1 U634 ( .A0(n24), .A1(n773), .B0(n772), .B1(n22), .Y(n640) );
  OAI22X1 U635 ( .A0(n24), .A1(n774), .B0(n773), .B1(n22), .Y(n641) );
  OAI22X1 U667 ( .A0(n18), .A1(n787), .B0(n786), .B1(n16), .Y(n653) );
  OAI22X1 U727 ( .A0(n6), .A1(n973), .B0(n827), .B1(n867), .Y(n563) );
  OAI22X1 U731 ( .A0(n6), .A1(n813), .B0(n812), .B1(n867), .Y(n678) );
  OAI22X1 U733 ( .A0(n6), .A1(n815), .B0(n814), .B1(n867), .Y(n680) );
  OAI22X1 U735 ( .A0(n6), .A1(n817), .B0(n816), .B1(n867), .Y(n682) );
  OAI22X1 U737 ( .A0(n6), .A1(n819), .B0(n818), .B1(n867), .Y(n684) );
  OAI22X1 U738 ( .A0(n6), .A1(n820), .B0(n819), .B1(n867), .Y(n685) );
  OAI22X1 U739 ( .A0(n6), .A1(n821), .B0(n820), .B1(n867), .Y(n686) );
  OAI22X1 U740 ( .A0(n6), .A1(n822), .B0(n821), .B1(n867), .Y(n687) );
  OAI22X1 U742 ( .A0(n6), .A1(n824), .B0(n823), .B1(n867), .Y(n689) );
  OAI22X1 U743 ( .A0(n6), .A1(n825), .B0(n824), .B1(n867), .Y(n690) );
  NAND2X4 U786 ( .A(n46), .B(n844), .Y(n48) );
  XNOR2X4 U788 ( .A(n1006), .B(a[14]), .Y(n46) );
  NAND2X4 U789 ( .A(n960), .B(n845), .Y(n42) );
  XNOR2X4 U791 ( .A(n1005), .B(a[12]), .Y(n40) );
  NAND2X4 U792 ( .A(n34), .B(n846), .Y(n36) );
  XNOR2X4 U794 ( .A(n1004), .B(a[10]), .Y(n34) );
  NAND2X4 U795 ( .A(n957), .B(n847), .Y(n30) );
  XNOR2X4 U797 ( .A(n1003), .B(a[8]), .Y(n28) );
  NAND2X4 U798 ( .A(n22), .B(n848), .Y(n24) );
  XNOR2X4 U800 ( .A(n1002), .B(a[6]), .Y(n22) );
  NAND2X4 U801 ( .A(n16), .B(n849), .Y(n18) );
  NAND2X4 U804 ( .A(n9), .B(n850), .Y(n12) );
  NAND2X4 U807 ( .A(n851), .B(n867), .Y(n6) );
  INVX2 U812 ( .A(n235), .Y(n954) );
  CLKINVX2 U813 ( .A(n1001), .Y(n969) );
  ADDFHX1 U814 ( .A(n668), .B(n523), .CI(n528), .CO(n518), .S(n519) );
  NOR2X2 U815 ( .A(n211), .B(n216), .Y(n209) );
  OAI21XL U816 ( .A0(n211), .A1(n219), .B0(n212), .Y(n210) );
  NOR2BXL U817 ( .AN(b[0]), .B(n16), .Y(n659) );
  OAI22XL U818 ( .A0(n18), .A1(n792), .B0(n791), .B1(n16), .Y(n658) );
  OAI22XL U819 ( .A0(n18), .A1(n788), .B0(n787), .B1(n16), .Y(n654) );
  OAI22XL U820 ( .A0(n18), .A1(n786), .B0(n785), .B1(n16), .Y(n652) );
  NOR2XL U821 ( .A(n6), .B(n812), .Y(n943) );
  NOR2XL U822 ( .A(n811), .B(n867), .Y(n944) );
  OR2X2 U823 ( .A(n943), .B(n944), .Y(n677) );
  INVX12 U824 ( .A(a[0]), .Y(n867) );
  OR2X4 U825 ( .A(n227), .B(n233), .Y(n945) );
  NAND2X4 U826 ( .A(n945), .B(n228), .Y(n222) );
  NAND2XL U827 ( .A(n437), .B(n450), .Y(n228) );
  AOI21X1 U828 ( .A0(n234), .A1(n221), .B0(n222), .Y(n220) );
  INVX2 U829 ( .A(n222), .Y(n224) );
  NAND2X4 U830 ( .A(n946), .B(n947), .Y(n948) );
  NAND2X4 U831 ( .A(n948), .B(n200), .Y(n194) );
  INVX3 U832 ( .A(n199), .Y(n946) );
  INVX4 U833 ( .A(n205), .Y(n947) );
  CLKINVX1 U834 ( .A(n194), .Y(n196) );
  OAI2BB1X4 U835 ( .A0N(n194), .A1N(n181), .B0(n989), .Y(n988) );
  AOI21XL U836 ( .A0(n51), .A1(n193), .B0(n194), .Y(n192) );
  OR2X4 U837 ( .A(n12), .B(n795), .Y(n949) );
  OR2X2 U838 ( .A(n794), .B(n9), .Y(n950) );
  NAND2X4 U839 ( .A(n949), .B(n950), .Y(n434) );
  XNOR2XL U840 ( .A(b[15]), .B(n1001), .Y(n794) );
  INVX3 U841 ( .A(n434), .Y(n435) );
  OR2X1 U842 ( .A(n18), .B(n789), .Y(n951) );
  OR2X1 U843 ( .A(n788), .B(n16), .Y(n952) );
  NAND2X2 U844 ( .A(n951), .B(n952), .Y(n655) );
  ADDFHX1 U845 ( .A(n669), .B(n655), .CI(n534), .CO(n526), .S(n527) );
  NAND2X2 U846 ( .A(n953), .B(n954), .Y(n955) );
  NAND2X4 U847 ( .A(n955), .B(n208), .Y(n51) );
  INVX2 U848 ( .A(n207), .Y(n953) );
  AOI21X1 U849 ( .A0(n51), .A1(n142), .B0(n143), .Y(n141) );
  AOI21X1 U850 ( .A0(n51), .A1(n155), .B0(n156), .Y(n154) );
  AOI21X1 U851 ( .A0(n51), .A1(n177), .B0(n988), .Y(n176) );
  XOR2X1 U852 ( .A(n51), .B(n987), .Y(product[19]) );
  ADDFX1 U853 ( .A(n604), .B(n646), .CI(n435), .CO(n432), .S(n433) );
  OAI21X2 U854 ( .A0(n242), .A1(n238), .B0(n239), .Y(n237) );
  AOI21X4 U855 ( .A0(n967), .A1(n251), .B0(n244), .Y(n242) );
  OAI22X1 U856 ( .A0(n12), .A1(n798), .B0(n797), .B1(n9), .Y(n663) );
  OAI22X1 U857 ( .A0(n6), .A1(n818), .B0(n817), .B1(n867), .Y(n683) );
  ADDFHX2 U858 ( .A(n635), .B(n964), .CI(n486), .CO(n470), .S(n471) );
  OAI22X2 U859 ( .A0(n24), .A1(n768), .B0(n767), .B1(n22), .Y(n635) );
  ADDFHX1 U860 ( .A(n647), .B(n577), .CI(n605), .CO(n444), .S(n445) );
  AOI21X1 U861 ( .A0(n51), .A1(n186), .B0(n187), .Y(n185) );
  AOI21X1 U862 ( .A0(n51), .A1(n168), .B0(n169), .Y(n167) );
  OAI22X1 U863 ( .A0(n12), .A1(n799), .B0(n798), .B1(n9), .Y(n664) );
  OAI22X1 U864 ( .A0(n36), .A1(n738), .B0(n737), .B1(n34), .Y(n607) );
  XNOR2X2 U865 ( .A(n167), .B(n980), .Y(product[24]) );
  INVX4 U866 ( .A(n28), .Y(n956) );
  CLKINVX3 U867 ( .A(n956), .Y(n957) );
  INVX16 U868 ( .A(n956), .Y(n958) );
  OAI22X1 U869 ( .A0(n18), .A1(n784), .B0(n783), .B1(n16), .Y(n650) );
  XNOR2XL U870 ( .A(b[4]), .B(n1002), .Y(n788) );
  XNOR2XL U871 ( .A(b[4]), .B(n1006), .Y(n720) );
  XNOR2XL U872 ( .A(b[4]), .B(n1004), .Y(n754) );
  INVX4 U873 ( .A(n40), .Y(n959) );
  CLKINVX4 U874 ( .A(n959), .Y(n960) );
  INVX2 U875 ( .A(n959), .Y(n961) );
  INVX1 U876 ( .A(n959), .Y(n962) );
  OAI22X2 U877 ( .A0(n30), .A1(n753), .B0(n752), .B1(n958), .Y(n621) );
  ADDFHX1 U878 ( .A(n622), .B(n594), .CI(n608), .CO(n482), .S(n483) );
  ADDFHX1 U879 ( .A(n638), .B(n624), .CI(n507), .CO(n502), .S(n503) );
  OAI22XL U880 ( .A0(n30), .A1(n756), .B0(n755), .B1(n958), .Y(n624) );
  XNOR2X1 U881 ( .A(b[3]), .B(n1004), .Y(n755) );
  XNOR2X1 U882 ( .A(b[3]), .B(n1005), .Y(n738) );
  OAI22X1 U883 ( .A0(n42), .A1(n869), .B0(n961), .B1(n725), .Y(n557) );
  ADDFHX2 U884 ( .A(n442), .B(n429), .CI(n440), .CO(n424), .S(n425) );
  ADDFHX2 U885 ( .A(n462), .B(n449), .CI(n460), .CO(n442), .S(n443) );
  ADDFHX1 U886 ( .A(n458), .B(n447), .CI(n445), .CO(n440), .S(n441) );
  ADDFHX1 U887 ( .A(n556), .B(n578), .CI(n592), .CO(n460), .S(n461) );
  OAI22XL U888 ( .A0(n48), .A1(n707), .B0(n706), .B1(n46), .Y(n578) );
  OAI22XL U889 ( .A0(n36), .A1(n729), .B0(n728), .B1(n34), .Y(n598) );
  OAI22XL U890 ( .A0(n36), .A1(n728), .B0(n727), .B1(n34), .Y(n597) );
  OAI22XL U891 ( .A0(n36), .A1(n727), .B0(n726), .B1(n34), .Y(n354) );
  OAI22XL U892 ( .A0(n36), .A1(n731), .B0(n730), .B1(n34), .Y(n600) );
  OAI22XL U893 ( .A0(n36), .A1(n732), .B0(n731), .B1(n34), .Y(n601) );
  OAI22XL U894 ( .A0(n36), .A1(n736), .B0(n735), .B1(n34), .Y(n605) );
  OAI22XL U895 ( .A0(n36), .A1(n734), .B0(n733), .B1(n34), .Y(n603) );
  OAI22XL U896 ( .A0(n36), .A1(n739), .B0(n738), .B1(n34), .Y(n608) );
  OAI22XL U897 ( .A0(n36), .A1(n733), .B0(n732), .B1(n34), .Y(n602) );
  OAI22XL U898 ( .A0(n36), .A1(n740), .B0(n739), .B1(n34), .Y(n609) );
  OAI22XL U899 ( .A0(n36), .A1(n735), .B0(n734), .B1(n34), .Y(n604) );
  ADDFHX1 U900 ( .A(n662), .B(n606), .CI(n620), .CO(n458), .S(n459) );
  XNOR2X1 U901 ( .A(b[13]), .B(n1002), .Y(n779) );
  XNOR2X1 U902 ( .A(b[13]), .B(n1003), .Y(n762) );
  XNOR2X1 U903 ( .A(b[13]), .B(n1000), .Y(n813) );
  XNOR2X1 U904 ( .A(b[13]), .B(n1001), .Y(n796) );
  INVX1 U905 ( .A(n607), .Y(n963) );
  INVX2 U906 ( .A(n963), .Y(n964) );
  ADDFHX1 U907 ( .A(n575), .B(n434), .CI(n660), .CO(n420), .S(n421) );
  ADDFHX1 U908 ( .A(n558), .B(n610), .CI(n666), .CO(n504), .S(n505) );
  OAI22XL U909 ( .A0(n36), .A1(n741), .B0(n740), .B1(n34), .Y(n610) );
  ADDFHX1 U910 ( .A(n621), .B(n663), .CI(n649), .CO(n472), .S(n473) );
  ADDFHX1 U911 ( .A(n557), .B(n664), .CI(n636), .CO(n484), .S(n485) );
  XOR2X2 U912 ( .A(a[14]), .B(n1007), .Y(n844) );
  XNOR2X1 U913 ( .A(b[9]), .B(n1003), .Y(n766) );
  XNOR2X1 U914 ( .A(b[9]), .B(n1002), .Y(n783) );
  XNOR2X1 U915 ( .A(b[9]), .B(n1005), .Y(n732) );
  XNOR2X1 U916 ( .A(b[9]), .B(n1001), .Y(n800) );
  XNOR2X1 U917 ( .A(b[10]), .B(n1001), .Y(n799) );
  XNOR2X1 U918 ( .A(b[10]), .B(n1003), .Y(n765) );
  XNOR2X1 U919 ( .A(b[15]), .B(n1002), .Y(n777) );
  XNOR2X1 U920 ( .A(b[12]), .B(n1001), .Y(n797) );
  XNOR2X1 U921 ( .A(b[12]), .B(n1002), .Y(n780) );
  XNOR2X1 U922 ( .A(b[12]), .B(n1003), .Y(n763) );
  AOI21XL U923 ( .A0(n51), .A1(n85), .B0(n86), .Y(product[31]) );
  AOI21XL U924 ( .A0(n51), .A1(n94), .B0(n95), .Y(n93) );
  AOI21XL U925 ( .A0(n51), .A1(n118), .B0(n119), .Y(n117) );
  AOI21XL U926 ( .A0(n51), .A1(n107), .B0(n108), .Y(n106) );
  XNOR2X1 U927 ( .A(b[11]), .B(n1001), .Y(n798) );
  XNOR2X1 U928 ( .A(b[11]), .B(n1000), .Y(n815) );
  XNOR2X1 U929 ( .A(b[11]), .B(n1002), .Y(n781) );
  XNOR2X1 U930 ( .A(b[11]), .B(n1003), .Y(n764) );
  BUFX8 U931 ( .A(a[7]), .Y(n1003) );
  BUFX8 U932 ( .A(a[9]), .Y(n1004) );
  BUFX8 U933 ( .A(a[11]), .Y(n1005) );
  OAI22XL U934 ( .A0(n24), .A1(n761), .B0(n760), .B1(n22), .Y(n386) );
  ADDFX1 U935 ( .A(n602), .B(n630), .CI(n409), .CO(n406), .S(n407) );
  ADDFX2 U936 ( .A(n585), .B(n599), .CI(n613), .CO(n374), .S(n375) );
  BUFX8 U937 ( .A(a[15]), .Y(n1007) );
  NAND2X2 U938 ( .A(n399), .B(n410), .Y(n205) );
  ADDFX2 U939 ( .A(n360), .B(n353), .CI(n358), .CO(n350), .S(n351) );
  ADDFX2 U940 ( .A(n581), .B(n352), .CI(n349), .CO(n346), .S(n347) );
  NOR2X2 U941 ( .A(n188), .B(n183), .Y(n181) );
  OAI22XL U942 ( .A0(n6), .A1(n823), .B0(n822), .B1(n867), .Y(n688) );
  ADDHXL U943 ( .A(n681), .B(n652), .CO(n506), .S(n507) );
  OAI21X1 U944 ( .A0(n298), .A1(n296), .B0(n297), .Y(n295) );
  NAND2BX1 U945 ( .AN(n1008), .B(n1007), .Y(n708) );
  XOR2X1 U946 ( .A(n262), .B(n73), .Y(product[11]) );
  NOR2X1 U947 ( .A(n489), .B(n498), .Y(n248) );
  ADDFX1 U948 ( .A(n571), .B(n386), .CI(n628), .CO(n376), .S(n377) );
  XOR2X1 U949 ( .A(n1005), .B(a[10]), .Y(n846) );
  NAND2X1 U950 ( .A(n477), .B(n488), .Y(n246) );
  INVX2 U951 ( .A(n248), .Y(n326) );
  ADDFX2 U952 ( .A(n584), .B(n570), .CI(n369), .CO(n366), .S(n367) );
  ADDFHX1 U953 ( .A(n441), .B(n452), .CI(n439), .CO(n436), .S(n437) );
  ADDFHX1 U954 ( .A(n427), .B(n438), .CI(n425), .CO(n422), .S(n423) );
  NAND2X2 U955 ( .A(n451), .B(n464), .Y(n233) );
  NOR2X2 U956 ( .A(n437), .B(n450), .Y(n227) );
  NAND2X2 U957 ( .A(n423), .B(n436), .Y(n219) );
  NOR2X1 U958 ( .A(n356), .B(n351), .Y(n148) );
  ADDFHX1 U959 ( .A(n367), .B(n365), .CI(n372), .CO(n362), .S(n363) );
  NAND2X1 U960 ( .A(n122), .B(n98), .Y(n96) );
  OAI21X1 U961 ( .A0(n158), .A1(n124), .B0(n125), .Y(n123) );
  NAND2X1 U962 ( .A(n356), .B(n351), .Y(n149) );
  NOR2X1 U963 ( .A(n370), .B(n363), .Y(n170) );
  CLKINVX2 U964 ( .A(n182), .Y(n989) );
  OAI21XL U965 ( .A0(n183), .A1(n191), .B0(n184), .Y(n182) );
  NOR2X1 U966 ( .A(n350), .B(n347), .Y(n137) );
  NOR2X1 U967 ( .A(n346), .B(n343), .Y(n128) );
  ADDHXL U968 ( .A(n689), .B(n562), .CO(n546), .S(n547) );
  NOR2X1 U969 ( .A(n24), .B(n775), .Y(n977) );
  NOR2X1 U970 ( .A(n774), .B(n22), .Y(n978) );
  OR2X2 U971 ( .A(n547), .B(n674), .Y(n996) );
  OAI21X1 U972 ( .A0(n304), .A1(n307), .B0(n305), .Y(n303) );
  ADDFX2 U973 ( .A(n559), .B(n626), .CI(n640), .CO(n520), .S(n521) );
  ADDFX2 U974 ( .A(n639), .B(n653), .CI(n667), .CO(n512), .S(n513) );
  ADDFX2 U975 ( .A(n637), .B(n665), .CI(n623), .CO(n494), .S(n495) );
  ADDFX2 U976 ( .A(n651), .B(n506), .CI(n497), .CO(n492), .S(n493) );
  NOR2X1 U977 ( .A(n690), .B(n675), .Y(n304) );
  AOI21X1 U978 ( .A0(n295), .A1(n994), .B0(n292), .Y(n290) );
  OR2X2 U979 ( .A(n531), .B(n536), .Y(n993) );
  NAND2X1 U980 ( .A(n509), .B(n516), .Y(n266) );
  ADDFX2 U981 ( .A(n521), .B(n526), .CI(n519), .CO(n516), .S(n517) );
  ADDFX2 U982 ( .A(n513), .B(n518), .CI(n511), .CO(n508), .S(n509) );
  ADDFHX1 U983 ( .A(n504), .B(n502), .CI(n495), .CO(n490), .S(n491) );
  ADDFX2 U984 ( .A(n487), .B(n496), .CI(n494), .CO(n480), .S(n481) );
  ADDFX2 U985 ( .A(n634), .B(n463), .CI(n474), .CO(n456), .S(n457) );
  ADDFX2 U986 ( .A(n632), .B(n576), .CI(n618), .CO(n430), .S(n431) );
  ADDFX2 U987 ( .A(n590), .B(n448), .CI(n446), .CO(n428), .S(n429) );
  XNOR2X1 U988 ( .A(n633), .B(n591), .Y(n449) );
  ADDFHX1 U989 ( .A(n485), .B(n483), .CI(n492), .CO(n478), .S(n479) );
  ADDFX2 U990 ( .A(n475), .B(n484), .CI(n473), .CO(n468), .S(n469) );
  ADDFX2 U991 ( .A(n472), .B(n470), .CI(n459), .CO(n454), .S(n455) );
  ADDFX2 U992 ( .A(n482), .B(n471), .CI(n480), .CO(n466), .S(n467) );
  ADDFX2 U993 ( .A(n645), .B(n589), .CI(n631), .CO(n418), .S(n419) );
  ADDFX2 U994 ( .A(n617), .B(n603), .CI(n432), .CO(n416), .S(n417) );
  ADDFX2 U995 ( .A(n629), .B(n587), .CI(n601), .CO(n394), .S(n395) );
  ADDFX2 U996 ( .A(n586), .B(n614), .CI(n387), .CO(n384), .S(n385) );
  OR2X1 U997 ( .A(n509), .B(n516), .Y(n992) );
  INVX2 U998 ( .A(n260), .Y(n327) );
  NOR2X1 U999 ( .A(n499), .B(n508), .Y(n260) );
  ADDFHX1 U1000 ( .A(n461), .B(n457), .CI(n468), .CO(n452), .S(n453) );
  ADDFX2 U1001 ( .A(n444), .B(n433), .CI(n431), .CO(n426), .S(n427) );
  ADDFHX1 U1002 ( .A(n456), .B(n443), .CI(n454), .CO(n438), .S(n439) );
  ADDFX2 U1003 ( .A(n430), .B(n421), .CI(n419), .CO(n414), .S(n415) );
  ADDFHX1 U1004 ( .A(n428), .B(n417), .CI(n426), .CO(n412), .S(n413) );
  ADDFX2 U1005 ( .A(n469), .B(n478), .CI(n467), .CO(n464), .S(n465) );
  XOR2X1 U1006 ( .A(n247), .B(n990), .Y(product[13]) );
  OAI21X1 U1007 ( .A0(n254), .A1(n248), .B0(n249), .Y(n247) );
  NAND2X1 U1008 ( .A(n324), .B(n239), .Y(n70) );
  ADDFX2 U1009 ( .A(n615), .B(n406), .CI(n404), .CO(n392), .S(n393) );
  ADDFX2 U1010 ( .A(n395), .B(n397), .CI(n393), .CO(n390), .S(n391) );
  ADDFX2 U1011 ( .A(n418), .B(n416), .CI(n414), .CO(n400), .S(n401) );
  ADDFX2 U1012 ( .A(n420), .B(n405), .CI(n407), .CO(n402), .S(n403) );
  ADDFX2 U1013 ( .A(n600), .B(n572), .CI(n396), .CO(n382), .S(n383) );
  ADDFX2 U1014 ( .A(n394), .B(n385), .CI(n383), .CO(n380), .S(n381) );
  ADDFX2 U1015 ( .A(n598), .B(n376), .CI(n374), .CO(n364), .S(n365) );
  ADDFX2 U1016 ( .A(n384), .B(n377), .CI(n375), .CO(n372), .S(n373) );
  ADDFX2 U1017 ( .A(n597), .B(n583), .CI(n366), .CO(n358), .S(n359) );
  ADDFX2 U1018 ( .A(n582), .B(n568), .CI(n355), .CO(n352), .S(n353) );
  NOR2X1 U1019 ( .A(n137), .B(n128), .Y(n126) );
  NOR2X2 U1020 ( .A(n465), .B(n476), .Y(n238) );
  INVX2 U1021 ( .A(n246), .Y(n244) );
  INVX2 U1022 ( .A(n249), .Y(n251) );
  NAND2X1 U1023 ( .A(n967), .B(n326), .Y(n241) );
  NAND2X1 U1024 ( .A(n465), .B(n476), .Y(n239) );
  NAND2X1 U1025 ( .A(n320), .B(n212), .Y(n66) );
  XOR2X1 U1026 ( .A(n229), .B(n68), .Y(product[16]) );
  NAND2X1 U1027 ( .A(n322), .B(n228), .Y(n68) );
  XOR2X1 U1028 ( .A(n220), .B(n67), .Y(product[17]) );
  NAND2X1 U1029 ( .A(n321), .B(n219), .Y(n67) );
  NOR2X1 U1030 ( .A(n227), .B(n232), .Y(n221) );
  NOR2X2 U1031 ( .A(n423), .B(n436), .Y(n216) );
  NOR2X2 U1032 ( .A(n411), .B(n422), .Y(n211) );
  AND2X1 U1033 ( .A(n319), .B(n205), .Y(n987) );
  XOR2X1 U1034 ( .A(n201), .B(n64), .Y(product[20]) );
  XOR2X1 U1035 ( .A(n192), .B(n63), .Y(product[21]) );
  XNOR2X1 U1036 ( .A(n154), .B(n981), .Y(product[25]) );
  NOR2X1 U1037 ( .A(n53), .B(n157), .Y(n155) );
  NOR2X1 U1038 ( .A(n53), .B(n170), .Y(n168) );
  NOR2X1 U1039 ( .A(n53), .B(n120), .Y(n118) );
  NOR2X1 U1040 ( .A(n53), .B(n109), .Y(n107) );
  XOR2X1 U1041 ( .A(n185), .B(n62), .Y(product[22]) );
  NOR2BX1 U1042 ( .AN(n193), .B(n188), .Y(n186) );
  XOR2X1 U1043 ( .A(n176), .B(n61), .Y(product[23]) );
  INVX2 U1044 ( .A(n53), .Y(n177) );
  XNOR2X1 U1045 ( .A(n141), .B(n984), .Y(product[26]) );
  XOR2X1 U1046 ( .A(n130), .B(n57), .Y(product[27]) );
  XNOR2X1 U1047 ( .A(n93), .B(n985), .Y(product[30]) );
  NOR2X1 U1048 ( .A(n53), .B(n87), .Y(n85) );
  NAND2X1 U1049 ( .A(n691), .B(n563), .Y(n307) );
  OAI22X1 U1050 ( .A0(n6), .A1(n826), .B0(n825), .B1(n867), .Y(n691) );
  INVX1 U1051 ( .A(n682), .Y(n965) );
  CLKINVX2 U1052 ( .A(n965), .Y(n966) );
  OAI21X1 U1053 ( .A0(n268), .A1(n256), .B0(n257), .Y(n255) );
  OR2X4 U1054 ( .A(n477), .B(n488), .Y(n967) );
  INVX2 U1055 ( .A(n988), .Y(n52) );
  OR2X1 U1056 ( .A(n691), .B(n563), .Y(n968) );
  NOR2X1 U1057 ( .A(n362), .B(n357), .Y(n165) );
  BUFX4 U1058 ( .A(a[3]), .Y(n1001) );
  BUFX4 U1059 ( .A(a[1]), .Y(n1000) );
  ADDFHX2 U1060 ( .A(n535), .B(n538), .CI(n533), .CO(n530), .S(n531) );
  NAND2X1 U1061 ( .A(n1001), .B(a[4]), .Y(n971) );
  NAND2X2 U1062 ( .A(n969), .B(n970), .Y(n972) );
  NAND2X4 U1063 ( .A(n971), .B(n972), .Y(n16) );
  INVX2 U1064 ( .A(a[4]), .Y(n970) );
  OAI22X1 U1065 ( .A0(n18), .A1(n780), .B0(n779), .B1(n16), .Y(n646) );
  OAI22XL U1066 ( .A0(n18), .A1(n791), .B0(n790), .B1(n16), .Y(n657) );
  OAI22XL U1067 ( .A0(n18), .A1(n785), .B0(n784), .B1(n16), .Y(n651) );
  OAI22XL U1068 ( .A0(n18), .A1(n778), .B0(n777), .B1(n16), .Y(n408) );
  OAI22XL U1069 ( .A0(n18), .A1(n873), .B0(n16), .B1(n793), .Y(n561) );
  OAI22XL U1070 ( .A0(n18), .A1(n782), .B0(n781), .B1(n16), .Y(n648) );
  OAI22XL U1071 ( .A0(n18), .A1(n783), .B0(n782), .B1(n16), .Y(n649) );
  OAI22XL U1072 ( .A0(n18), .A1(n779), .B0(n778), .B1(n16), .Y(n645) );
  NAND2X1 U1073 ( .A(n1000), .B(a[2]), .Y(n975) );
  NAND2X2 U1074 ( .A(n973), .B(n974), .Y(n976) );
  NAND2X4 U1075 ( .A(n975), .B(n976), .Y(n9) );
  CLKINVXL U1076 ( .A(n1000), .Y(n973) );
  INVX2 U1077 ( .A(a[2]), .Y(n974) );
  OAI22XL U1078 ( .A0(n12), .A1(n807), .B0(n806), .B1(n9), .Y(n672) );
  OAI22XL U1079 ( .A0(n12), .A1(n805), .B0(n804), .B1(n9), .Y(n670) );
  OAI22XL U1080 ( .A0(n12), .A1(n797), .B0(n796), .B1(n9), .Y(n662) );
  OAI22XL U1081 ( .A0(n12), .A1(n806), .B0(n805), .B1(n9), .Y(n671) );
  OAI22XL U1082 ( .A0(n12), .A1(n801), .B0(n800), .B1(n9), .Y(n666) );
  OAI22XL U1083 ( .A0(n12), .A1(n809), .B0(n808), .B1(n9), .Y(n674) );
  OAI22XL U1084 ( .A0(n12), .A1(n808), .B0(n807), .B1(n9), .Y(n673) );
  OAI22XL U1085 ( .A0(n12), .A1(n969), .B0(n9), .B1(n810), .Y(n562) );
  OAI22XL U1086 ( .A0(n12), .A1(n804), .B0(n803), .B1(n9), .Y(n669) );
  OAI22XL U1087 ( .A0(n12), .A1(n796), .B0(n795), .B1(n9), .Y(n661) );
  OAI22XL U1088 ( .A0(n12), .A1(n803), .B0(n802), .B1(n9), .Y(n668) );
  OAI22XL U1089 ( .A0(n12), .A1(n802), .B0(n801), .B1(n9), .Y(n667) );
  CLKINVXL U1090 ( .A(n1009), .Y(n1008) );
  XNOR2XL U1091 ( .A(b[1]), .B(n1003), .Y(n774) );
  OR2X1 U1092 ( .A(n977), .B(n978), .Y(n642) );
  XNOR2XL U1093 ( .A(b[0]), .B(n1003), .Y(n775) );
  AOI2BB1X1 U1094 ( .A0N(n165), .A1N(n171), .B0(n164), .Y(n158) );
  CLKINVXL U1095 ( .A(n232), .Y(n323) );
  NAND2X2 U1096 ( .A(n411), .B(n422), .Y(n212) );
  NAND2X1 U1097 ( .A(n690), .B(n675), .Y(n305) );
  NAND2BXL U1098 ( .AN(n1008), .B(n1005), .Y(n742) );
  INVX1 U1099 ( .A(n268), .Y(n267) );
  AOI21X2 U1100 ( .A0(n209), .A1(n222), .B0(n210), .Y(n208) );
  OAI21XL U1101 ( .A0(n268), .A1(n256), .B0(n257), .Y(n986) );
  AOI21XL U1102 ( .A0(n51), .A1(n319), .B0(n203), .Y(n201) );
  XOR2X1 U1103 ( .A(n234), .B(n979), .Y(product[15]) );
  AND2X1 U1104 ( .A(n323), .B(n233), .Y(n979) );
  OAI21XL U1105 ( .A0(n254), .A1(n241), .B0(n242), .Y(n240) );
  CLKINVXL U1106 ( .A(n238), .Y(n324) );
  INVX2 U1107 ( .A(n204), .Y(n319) );
  INVX2 U1108 ( .A(n157), .Y(n159) );
  NOR2X1 U1109 ( .A(n157), .B(n124), .Y(n122) );
  AOI21X1 U1110 ( .A0(n267), .A1(n992), .B0(n264), .Y(n262) );
  INVX2 U1111 ( .A(n266), .Y(n264) );
  NAND2XL U1112 ( .A(n315), .B(n171), .Y(n61) );
  NAND2X1 U1113 ( .A(n159), .B(n135), .Y(n133) );
  INVX2 U1114 ( .A(n170), .Y(n315) );
  NAND2X1 U1115 ( .A(n313), .B(n126), .Y(n124) );
  INVX2 U1116 ( .A(n148), .Y(n313) );
  INVX1 U1117 ( .A(n294), .Y(n292) );
  INVX1 U1118 ( .A(n288), .Y(n286) );
  NAND2X1 U1119 ( .A(n499), .B(n508), .Y(n261) );
  AOI21XL U1120 ( .A0(n51), .A1(n131), .B0(n132), .Y(n130) );
  NAND2X2 U1121 ( .A(n379), .B(n388), .Y(n191) );
  ADDFHX1 U1122 ( .A(n560), .B(n642), .CI(n670), .CO(n532), .S(n533) );
  ADDHX1 U1123 ( .A(n677), .B(n648), .CO(n462), .S(n463) );
  OR2X1 U1124 ( .A(n633), .B(n591), .Y(n448) );
  OAI22XL U1125 ( .A0(n42), .A1(n724), .B0(n723), .B1(n962), .Y(n594) );
  ADDHXL U1126 ( .A(n679), .B(n650), .CO(n486), .S(n487) );
  ADDFX2 U1127 ( .A(n566), .B(n345), .CI(n348), .CO(n342), .S(n343) );
  XOR2X1 U1128 ( .A(n1004), .B(a[8]), .Y(n847) );
  XNOR2XL U1129 ( .A(b[4]), .B(n1003), .Y(n771) );
  XOR2X1 U1130 ( .A(n1006), .B(a[12]), .Y(n845) );
  XNOR2XL U1131 ( .A(b[3]), .B(n1006), .Y(n721) );
  XNOR2XL U1132 ( .A(b[2]), .B(n1006), .Y(n722) );
  XNOR2XL U1133 ( .A(b[8]), .B(n1006), .Y(n716) );
  XNOR2XL U1134 ( .A(b[10]), .B(n1006), .Y(n714) );
  XNOR2XL U1135 ( .A(b[9]), .B(n1006), .Y(n715) );
  XNOR2XL U1136 ( .A(b[10]), .B(n1005), .Y(n731) );
  XNOR2XL U1137 ( .A(b[10]), .B(n1007), .Y(n697) );
  XNOR2XL U1138 ( .A(b[12]), .B(n1007), .Y(n695) );
  XNOR2XL U1139 ( .A(b[14]), .B(n1007), .Y(n693) );
  XNOR2X1 U1140 ( .A(n240), .B(n70), .Y(product[14]) );
  XOR2X1 U1141 ( .A(n213), .B(n66), .Y(product[18]) );
  AOI21XL U1142 ( .A0(n214), .A1(n234), .B0(n215), .Y(n213) );
  AOI21XL U1143 ( .A0(n234), .A1(n323), .B0(n231), .Y(n229) );
  NAND2BX1 U1144 ( .AN(n199), .B(n200), .Y(n64) );
  OAI21XL U1145 ( .A0(n52), .A1(n157), .B0(n158), .Y(n156) );
  NAND2X1 U1146 ( .A(n159), .B(n313), .Y(n144) );
  XOR2X1 U1147 ( .A(n254), .B(n72), .Y(product[12]) );
  NAND2XL U1148 ( .A(n329), .B(n272), .Y(n75) );
  OAI21XL U1149 ( .A0(n276), .A1(n274), .B0(n275), .Y(n273) );
  CLKINVXL U1150 ( .A(n271), .Y(n329) );
  CLKINVXL U1151 ( .A(n277), .Y(n276) );
  XOR2X1 U1152 ( .A(n276), .B(n76), .Y(product[8]) );
  NAND2XL U1153 ( .A(n330), .B(n275), .Y(n76) );
  CLKINVXL U1154 ( .A(n274), .Y(n330) );
  NAND2BX1 U1155 ( .AN(n183), .B(n184), .Y(n62) );
  NAND2BX1 U1156 ( .AN(n188), .B(n191), .Y(n63) );
  AND2X1 U1157 ( .A(n314), .B(n166), .Y(n980) );
  AND2X1 U1158 ( .A(n313), .B(n149), .Y(n981) );
  NAND2X1 U1159 ( .A(n389), .B(n398), .Y(n200) );
  OAI21XL U1160 ( .A0(n52), .A1(n96), .B0(n97), .Y(n95) );
  INVX2 U1161 ( .A(n149), .Y(n151) );
  NAND2XL U1162 ( .A(n122), .B(n89), .Y(n87) );
  XOR2X1 U1163 ( .A(n80), .B(n298), .Y(product[4]) );
  NAND2XL U1164 ( .A(n334), .B(n297), .Y(n80) );
  CLKINVXL U1165 ( .A(n296), .Y(n334) );
  XOR2X1 U1166 ( .A(n284), .B(n77), .Y(product[7]) );
  AOI21XL U1167 ( .A0(n289), .A1(n995), .B0(n286), .Y(n284) );
  XOR2X1 U1168 ( .A(n982), .B(n289), .Y(product[6]) );
  AND2X1 U1169 ( .A(n995), .B(n288), .Y(n982) );
  XOR2XL U1170 ( .A(n983), .B(n295), .Y(product[5]) );
  AND2X1 U1171 ( .A(n994), .B(n294), .Y(n983) );
  AND2X1 U1172 ( .A(n312), .B(n140), .Y(n984) );
  XOR2XL U1173 ( .A(n82), .B(n307), .Y(product[2]) );
  CLKINVXL U1174 ( .A(n304), .Y(n336) );
  NAND2BX1 U1175 ( .AN(n128), .B(n129), .Y(n57) );
  AND2X1 U1176 ( .A(n308), .B(n92), .Y(n985) );
  XNOR2XL U1177 ( .A(n81), .B(n303), .Y(product[3]) );
  NAND2XL U1178 ( .A(n996), .B(n302), .Y(n81) );
  XOR2X1 U1179 ( .A(n106), .B(n55), .Y(product[29]) );
  XOR2X1 U1180 ( .A(n117), .B(n56), .Y(product[28]) );
  INVX2 U1181 ( .A(n165), .Y(n314) );
  AOI21XL U1182 ( .A0(n126), .A1(n151), .B0(n127), .Y(n125) );
  NAND2XL U1183 ( .A(n362), .B(n357), .Y(n166) );
  NAND2XL U1184 ( .A(n122), .B(n999), .Y(n109) );
  ADDFHX1 U1185 ( .A(n514), .B(n512), .CI(n505), .CO(n500), .S(n501) );
  ADDFHX1 U1186 ( .A(n522), .B(n515), .CI(n520), .CO(n510), .S(n511) );
  NAND2XL U1187 ( .A(n531), .B(n536), .Y(n283) );
  CMPR32X1 U1188 ( .A(n529), .B(n532), .C(n527), .CO(n524), .S(n525) );
  AND2X1 U1189 ( .A(n968), .B(n307), .Y(product[1]) );
  ADDHX1 U1190 ( .A(n683), .B(n654), .CO(n522), .S(n523) );
  XNOR2XL U1191 ( .A(b[0]), .B(n1002), .Y(n792) );
  CLKINVXL U1192 ( .A(n1002), .Y(n873) );
  CMPR32X1 U1193 ( .A(n672), .B(n561), .C(n543), .CO(n540), .S(n541) );
  ADDFHX1 U1194 ( .A(n643), .B(n686), .CI(n657), .CO(n538), .S(n539) );
  ADDFHX1 U1195 ( .A(n659), .B(n688), .CI(n673), .CO(n544), .S(n545) );
  ADDFX2 U1196 ( .A(n671), .B(n542), .CI(n539), .CO(n536), .S(n537) );
  OAI22XL U1197 ( .A0(n30), .A1(n871), .B0(n958), .B1(n759), .Y(n559) );
  OAI22XL U1198 ( .A0(n18), .A1(n790), .B0(n789), .B1(n16), .Y(n656) );
  OAI22XL U1199 ( .A0(n6), .A1(n816), .B0(n815), .B1(n867), .Y(n681) );
  NAND2BXL U1200 ( .AN(b[0]), .B(n1000), .Y(n827) );
  NAND2BXL U1201 ( .AN(n1008), .B(n1003), .Y(n776) );
  OAI22XL U1202 ( .A0(n42), .A1(n720), .B0(n719), .B1(n962), .Y(n590) );
  OAI22XL U1203 ( .A0(n36), .A1(n737), .B0(n736), .B1(n34), .Y(n606) );
  OAI22XL U1204 ( .A0(n12), .A1(n800), .B0(n799), .B1(n9), .Y(n665) );
  OAI22XL U1205 ( .A0(n6), .A1(n814), .B0(n813), .B1(n867), .Y(n679) );
  OAI22XL U1206 ( .A0(n18), .A1(n781), .B0(n780), .B1(n16), .Y(n647) );
  CLKINVXL U1207 ( .A(n1003), .Y(n872) );
  NAND2BXL U1208 ( .AN(n1008), .B(n1001), .Y(n810) );
  NAND2BXL U1209 ( .AN(n1008), .B(n1002), .Y(n793) );
  CLKINVXL U1210 ( .A(n1005), .Y(n870) );
  CLKINVXL U1211 ( .A(n794), .Y(n554) );
  CLKINVXL U1212 ( .A(n1004), .Y(n871) );
  OAI22XL U1213 ( .A0(n24), .A1(n765), .B0(n764), .B1(n22), .Y(n632) );
  OAI22XL U1214 ( .A0(n48), .A1(n701), .B0(n700), .B1(n46), .Y(n572) );
  OAI22XL U1215 ( .A0(n42), .A1(n719), .B0(n718), .B1(n961), .Y(n589) );
  CLKINVXL U1216 ( .A(n1006), .Y(n869) );
  OAI22XL U1217 ( .A0(n42), .A1(n717), .B0(n716), .B1(n961), .Y(n587) );
  INVX1 U1218 ( .A(n386), .Y(n387) );
  OAI22XL U1219 ( .A0(n42), .A1(n716), .B0(n715), .B1(n961), .Y(n586) );
  CLKINVXL U1220 ( .A(n760), .Y(n552) );
  INVXL U1221 ( .A(n368), .Y(n369) );
  OAI22XL U1222 ( .A0(n42), .A1(n714), .B0(n713), .B1(n961), .Y(n584) );
  OAI22XL U1223 ( .A0(n36), .A1(n730), .B0(n729), .B1(n34), .Y(n599) );
  OAI22XL U1224 ( .A0(n48), .A1(n697), .B0(n696), .B1(n46), .Y(n568) );
  XOR2X2 U1225 ( .A(n1000), .B(a[0]), .Y(n851) );
  XNOR2X1 U1226 ( .A(b[4]), .B(n1005), .Y(n737) );
  XNOR2X1 U1227 ( .A(b[1]), .B(n1006), .Y(n723) );
  XNOR2X1 U1228 ( .A(b[5]), .B(n1005), .Y(n736) );
  XNOR2X1 U1229 ( .A(b[4]), .B(n1007), .Y(n703) );
  XNOR2X1 U1230 ( .A(b[2]), .B(n1007), .Y(n705) );
  XNOR2X1 U1231 ( .A(b[1]), .B(n1007), .Y(n706) );
  XNOR2X1 U1232 ( .A(b[6]), .B(n1005), .Y(n735) );
  XNOR2XL U1233 ( .A(b[15]), .B(n1000), .Y(n811) );
  XNOR2X1 U1234 ( .A(b[3]), .B(n1007), .Y(n704) );
  XNOR2X1 U1235 ( .A(b[5]), .B(n1007), .Y(n702) );
  XNOR2X1 U1236 ( .A(b[6]), .B(n1007), .Y(n701) );
  XNOR2X1 U1237 ( .A(b[7]), .B(n1006), .Y(n717) );
  XNOR2X1 U1238 ( .A(b[5]), .B(n1006), .Y(n719) );
  XNOR2X1 U1239 ( .A(b[6]), .B(n1006), .Y(n718) );
  XNOR2X1 U1240 ( .A(b[8]), .B(n1007), .Y(n699) );
  XNOR2X1 U1241 ( .A(b[7]), .B(n1007), .Y(n700) );
  XNOR2X1 U1242 ( .A(b[9]), .B(n1007), .Y(n698) );
  XNOR2XL U1243 ( .A(b[13]), .B(n1007), .Y(n694) );
  XNOR2XL U1244 ( .A(b[15]), .B(n1007), .Y(n692) );
  NOR2XL U1245 ( .A(n53), .B(n96), .Y(n94) );
  INVX2 U1246 ( .A(n122), .Y(n120) );
  NOR2X1 U1247 ( .A(n53), .B(n144), .Y(n142) );
  CLKINVXL U1248 ( .A(n227), .Y(n322) );
  CLKINVXL U1249 ( .A(n216), .Y(n321) );
  INVX2 U1250 ( .A(n986), .Y(n254) );
  CLKINVXL U1251 ( .A(n211), .Y(n320) );
  NOR2BXL U1252 ( .AN(n221), .B(n216), .Y(n214) );
  OAI21XL U1253 ( .A0(n224), .A1(n216), .B0(n219), .Y(n215) );
  INVX2 U1254 ( .A(n158), .Y(n160) );
  OAI21XL U1255 ( .A0(n52), .A1(n144), .B0(n145), .Y(n143) );
  NOR2X1 U1256 ( .A(n53), .B(n133), .Y(n131) );
  CLKINVXL U1257 ( .A(n233), .Y(n231) );
  CLKINVXL U1258 ( .A(n205), .Y(n203) );
  INVX2 U1259 ( .A(n166), .Y(n164) );
  INVX2 U1260 ( .A(n101), .Y(n99) );
  NAND2X1 U1261 ( .A(n327), .B(n992), .Y(n256) );
  INVX2 U1262 ( .A(n261), .Y(n259) );
  AOI21X1 U1263 ( .A0(n269), .A1(n277), .B0(n270), .Y(n268) );
  OAI21X1 U1264 ( .A0(n271), .A1(n275), .B0(n272), .Y(n270) );
  NOR2X1 U1265 ( .A(n271), .B(n274), .Y(n269) );
  AND2X1 U1266 ( .A(n967), .B(n246), .Y(n990) );
  NAND2X1 U1267 ( .A(n327), .B(n261), .Y(n73) );
  NAND2X1 U1268 ( .A(n315), .B(n314), .Y(n157) );
  NAND2XL U1269 ( .A(n326), .B(n249), .Y(n72) );
  XNOR2X1 U1270 ( .A(n273), .B(n75), .Y(product[9]) );
  OAI21XL U1271 ( .A0(n52), .A1(n87), .B0(n88), .Y(n86) );
  INVX2 U1272 ( .A(n290), .Y(n289) );
  OAI21XL U1273 ( .A0(n52), .A1(n170), .B0(n171), .Y(n169) );
  NOR2X2 U1274 ( .A(n451), .B(n464), .Y(n232) );
  OAI21XL U1275 ( .A0(n52), .A1(n120), .B0(n121), .Y(n119) );
  CLKINVXL U1276 ( .A(n123), .Y(n121) );
  XOR2X1 U1277 ( .A(n267), .B(n991), .Y(product[10]) );
  AND2X1 U1278 ( .A(n992), .B(n266), .Y(n991) );
  OAI21XL U1279 ( .A0(n196), .A1(n188), .B0(n191), .Y(n187) );
  INVX2 U1280 ( .A(n100), .Y(n98) );
  OAI21XL U1281 ( .A0(n140), .A1(n128), .B0(n129), .Y(n127) );
  INVX2 U1282 ( .A(n91), .Y(n308) );
  NOR2X1 U1283 ( .A(n517), .B(n524), .Y(n271) );
  NOR2X1 U1284 ( .A(n525), .B(n530), .Y(n274) );
  OAI21XL U1285 ( .A0(n52), .A1(n109), .B0(n110), .Y(n108) );
  NAND2X1 U1286 ( .A(n998), .B(n105), .Y(n55) );
  OAI21X1 U1287 ( .A0(n278), .A1(n290), .B0(n279), .Y(n277) );
  AOI21X1 U1288 ( .A0(n993), .A1(n286), .B0(n281), .Y(n279) );
  NAND2X1 U1289 ( .A(n993), .B(n995), .Y(n278) );
  INVX2 U1290 ( .A(n283), .Y(n281) );
  OAI21X1 U1291 ( .A0(n101), .A1(n91), .B0(n92), .Y(n90) );
  NAND2X1 U1292 ( .A(n517), .B(n524), .Y(n272) );
  AOI21X2 U1293 ( .A0(n996), .A1(n303), .B0(n300), .Y(n298) );
  INVX2 U1294 ( .A(n302), .Y(n300) );
  NAND2X2 U1295 ( .A(n370), .B(n363), .Y(n171) );
  NAND2X1 U1296 ( .A(n999), .B(n116), .Y(n56) );
  NAND2X1 U1297 ( .A(n525), .B(n530), .Y(n275) );
  OAI21XL U1298 ( .A0(n52), .A1(n133), .B0(n134), .Y(n132) );
  OAI21XL U1299 ( .A0(n149), .A1(n137), .B0(n140), .Y(n136) );
  NAND2X1 U1300 ( .A(n993), .B(n283), .Y(n77) );
  NAND2X1 U1301 ( .A(n336), .B(n305), .Y(n82) );
  CLKINVXL U1302 ( .A(n137), .Y(n312) );
  NAND2X2 U1303 ( .A(n378), .B(n371), .Y(n184) );
  NOR2X1 U1304 ( .A(n148), .B(n137), .Y(n135) );
  INVX2 U1305 ( .A(n105), .Y(n103) );
  INVX2 U1306 ( .A(n116), .Y(n114) );
  NAND2X1 U1307 ( .A(n999), .B(n998), .Y(n100) );
  NOR2X1 U1308 ( .A(n100), .B(n91), .Y(n89) );
  OR2X1 U1309 ( .A(n541), .B(n544), .Y(n994) );
  OR2X1 U1310 ( .A(n537), .B(n540), .Y(n995) );
  NOR2X1 U1311 ( .A(n545), .B(n546), .Y(n296) );
  NAND2X1 U1312 ( .A(n541), .B(n544), .Y(n294) );
  NAND2X1 U1313 ( .A(n537), .B(n540), .Y(n288) );
  NAND2X1 U1314 ( .A(n547), .B(n674), .Y(n302) );
  NAND2X1 U1315 ( .A(n350), .B(n347), .Y(n140) );
  NAND2X1 U1316 ( .A(n545), .B(n546), .Y(n297) );
  NAND2XL U1317 ( .A(n346), .B(n343), .Y(n129) );
  NAND2X1 U1318 ( .A(n342), .B(n341), .Y(n116) );
  OR2X1 U1319 ( .A(n340), .B(n339), .Y(n998) );
  OR2X1 U1320 ( .A(n342), .B(n341), .Y(n999) );
  INVX2 U1321 ( .A(n338), .Y(n339) );
  NAND2X1 U1322 ( .A(n340), .B(n339), .Y(n105) );
  NOR2X1 U1323 ( .A(n564), .B(n338), .Y(n91) );
  NAND2X1 U1324 ( .A(n564), .B(n338), .Y(n92) );
  INVX2 U1325 ( .A(b[0]), .Y(n1009) );
  ADDFHX1 U1326 ( .A(n619), .B(n661), .CI(n676), .CO(n446), .S(n447) );
  OAI2BB1X1 U1327 ( .A0N(n867), .A1N(n6), .B0(n555), .Y(n676) );
  OAI22XL U1328 ( .A0(n36), .A1(n870), .B0(n34), .B1(n742), .Y(n558) );
  OAI2BB1X1 U1329 ( .A0N(n9), .A1N(n12), .B0(n554), .Y(n660) );
  ADDFX1 U1330 ( .A(n354), .B(n567), .CI(n596), .CO(n348), .S(n349) );
  OAI2BB1X1 U1331 ( .A0N(n34), .A1N(n36), .B0(n550), .Y(n596) );
  INVX2 U1332 ( .A(n726), .Y(n550) );
  NAND2BX1 U1333 ( .AN(n1008), .B(n1006), .Y(n725) );
  ADDFHX1 U1334 ( .A(n595), .B(n680), .CI(n609), .CO(n496), .S(n497) );
  ADDFHX1 U1335 ( .A(n627), .B(n684), .CI(n641), .CO(n528), .S(n529) );
  ADDHXL U1336 ( .A(n685), .B(n656), .CO(n534), .S(n535) );
  ADDFHX1 U1337 ( .A(n611), .B(n966), .CI(n625), .CO(n514), .S(n515) );
  XNOR2X1 U1338 ( .A(b[0]), .B(n1004), .Y(n758) );
  ADDFX1 U1339 ( .A(n579), .B(n678), .CI(n593), .CO(n474), .S(n475) );
  XNOR2X1 U1340 ( .A(b[0]), .B(n1006), .Y(n724) );
  INVX2 U1341 ( .A(n408), .Y(n409) );
  OAI22XL U1342 ( .A0(n24), .A1(n872), .B0(n22), .B1(n776), .Y(n560) );
  ADDFX1 U1343 ( .A(n569), .B(n368), .CI(n612), .CO(n360), .S(n361) );
  OAI2BB1X1 U1344 ( .A0N(n958), .A1N(n30), .B0(n551), .Y(n612) );
  INVX2 U1345 ( .A(n743), .Y(n551) );
  OAI2BB1X1 U1346 ( .A0N(n22), .A1N(n24), .B0(n552), .Y(n628) );
  XNOR2X1 U1347 ( .A(b[0]), .B(n1007), .Y(n707) );
  ADDFHX1 U1348 ( .A(n573), .B(n408), .CI(n644), .CO(n396), .S(n397) );
  OAI2BB1X1 U1349 ( .A0N(n16), .A1N(n18), .B0(n553), .Y(n644) );
  INVX2 U1350 ( .A(n777), .Y(n553) );
  ADDFHX1 U1351 ( .A(n574), .B(n588), .CI(n616), .CO(n404), .S(n405) );
  ADDHXL U1352 ( .A(n687), .B(n658), .CO(n542), .S(n543) );
  INVX2 U1353 ( .A(n344), .Y(n345) );
  CLKINVXL U1354 ( .A(n354), .Y(n355) );
  XNOR2X1 U1355 ( .A(b[0]), .B(n1000), .Y(n826) );
  ADDFX2 U1356 ( .A(n344), .B(n565), .CI(n580), .CO(n340), .S(n341) );
  OAI2BB1X1 U1357 ( .A0N(n961), .A1N(n42), .B0(n549), .Y(n580) );
  INVX2 U1358 ( .A(n709), .Y(n549) );
  INVX2 U1359 ( .A(n1007), .Y(n868) );
  INVX2 U1360 ( .A(n811), .Y(n555) );
  OAI2BB1X1 U1361 ( .A0N(n46), .A1N(n48), .B0(n548), .Y(n564) );
  INVX2 U1362 ( .A(n692), .Y(n548) );
  XOR2X1 U1363 ( .A(n1001), .B(a[2]), .Y(n850) );
  XOR2X1 U1364 ( .A(n1003), .B(a[6]), .Y(n848) );
  BUFX12 U1365 ( .A(a[5]), .Y(n1002) );
  XOR2X1 U1366 ( .A(n1002), .B(a[4]), .Y(n849) );
  BUFX12 U1367 ( .A(a[13]), .Y(n1006) );
  XNOR2XL U1368 ( .A(b[9]), .B(n1000), .Y(n817) );
  XNOR2XL U1369 ( .A(b[10]), .B(n1000), .Y(n816) );
  XNOR2XL U1370 ( .A(b[12]), .B(n1000), .Y(n814) );
  XNOR2XL U1371 ( .A(b[8]), .B(n1000), .Y(n818) );
  XNOR2XL U1372 ( .A(b[14]), .B(n1000), .Y(n812) );
  XNOR2XL U1373 ( .A(b[7]), .B(n1000), .Y(n819) );
  XNOR2XL U1374 ( .A(b[6]), .B(n1000), .Y(n820) );
  XNOR2XL U1375 ( .A(b[5]), .B(n1000), .Y(n821) );
  XNOR2X1 U1376 ( .A(b[4]), .B(n1000), .Y(n822) );
  XNOR2XL U1377 ( .A(b[15]), .B(n1004), .Y(n743) );
  XNOR2XL U1378 ( .A(b[14]), .B(n1001), .Y(n795) );
  XNOR2XL U1379 ( .A(b[15]), .B(n1005), .Y(n726) );
  XNOR2XL U1380 ( .A(b[7]), .B(n1002), .Y(n785) );
  XNOR2XL U1381 ( .A(b[14]), .B(n1004), .Y(n744) );
  XNOR2XL U1382 ( .A(b[6]), .B(n1004), .Y(n752) );
  XNOR2XL U1383 ( .A(b[5]), .B(n1002), .Y(n787) );
  XNOR2XL U1384 ( .A(b[3]), .B(n1002), .Y(n789) );
  XNOR2XL U1385 ( .A(b[6]), .B(n1002), .Y(n786) );
  XNOR2XL U1386 ( .A(b[8]), .B(n1004), .Y(n750) );
  XNOR2XL U1387 ( .A(b[8]), .B(n1002), .Y(n784) );
  XNOR2XL U1388 ( .A(b[3]), .B(n1000), .Y(n823) );
  XNOR2XL U1389 ( .A(b[14]), .B(n1005), .Y(n727) );
  XNOR2XL U1390 ( .A(b[5]), .B(n1004), .Y(n753) );
  XNOR2XL U1391 ( .A(b[7]), .B(n1005), .Y(n734) );
  XNOR2XL U1392 ( .A(b[10]), .B(n1002), .Y(n782) );
  XNOR2XL U1393 ( .A(b[15]), .B(n1003), .Y(n760) );
  XNOR2XL U1394 ( .A(b[1]), .B(n1000), .Y(n825) );
  XNOR2XL U1395 ( .A(b[2]), .B(n1002), .Y(n790) );
  XNOR2XL U1396 ( .A(b[1]), .B(n1005), .Y(n740) );
  XNOR2XL U1397 ( .A(b[1]), .B(n1004), .Y(n757) );
  XNOR2XL U1398 ( .A(b[7]), .B(n1004), .Y(n751) );
  XNOR2XL U1399 ( .A(b[2]), .B(n1000), .Y(n824) );
  XNOR2XL U1400 ( .A(b[3]), .B(n1003), .Y(n772) );
  XNOR2XL U1401 ( .A(b[8]), .B(n1005), .Y(n733) );
  XNOR2XL U1402 ( .A(b[6]), .B(n1003), .Y(n769) );
  XNOR2XL U1403 ( .A(b[14]), .B(n1002), .Y(n778) );
  XNOR2XL U1404 ( .A(b[1]), .B(n1002), .Y(n791) );
  XNOR2XL U1405 ( .A(b[8]), .B(n1003), .Y(n767) );
  XNOR2XL U1406 ( .A(b[14]), .B(n1003), .Y(n761) );
  XNOR2XL U1407 ( .A(b[13]), .B(n1004), .Y(n745) );
  XNOR2XL U1408 ( .A(b[2]), .B(n1005), .Y(n739) );
  XNOR2XL U1409 ( .A(b[2]), .B(n1004), .Y(n756) );
  XNOR2XL U1410 ( .A(b[5]), .B(n1003), .Y(n770) );
  XNOR2XL U1411 ( .A(b[12]), .B(n1005), .Y(n729) );
  XNOR2XL U1412 ( .A(b[7]), .B(n1003), .Y(n768) );
  XNOR2XL U1413 ( .A(b[6]), .B(n1001), .Y(n803) );
  XNOR2XL U1414 ( .A(b[12]), .B(n1004), .Y(n746) );
  XNOR2XL U1415 ( .A(b[11]), .B(n1006), .Y(n713) );
  XNOR2XL U1416 ( .A(b[2]), .B(n1003), .Y(n773) );
  XNOR2XL U1417 ( .A(b[11]), .B(n1005), .Y(n730) );
  XNOR2XL U1418 ( .A(b[5]), .B(n1001), .Y(n804) );
  XNOR2X1 U1419 ( .A(b[11]), .B(n1007), .Y(n696) );
  XNOR2XL U1420 ( .A(b[8]), .B(n1001), .Y(n801) );
  XNOR2XL U1421 ( .A(b[7]), .B(n1001), .Y(n802) );
  XNOR2XL U1422 ( .A(b[3]), .B(n1001), .Y(n806) );
  XNOR2XL U1423 ( .A(b[2]), .B(n1001), .Y(n807) );
  XNOR2XL U1424 ( .A(b[13]), .B(n1006), .Y(n711) );
  XNOR2X1 U1425 ( .A(b[4]), .B(n1001), .Y(n805) );
  XNOR2XL U1426 ( .A(b[1]), .B(n1001), .Y(n808) );
  XNOR2XL U1427 ( .A(b[9]), .B(n1004), .Y(n749) );
  XNOR2XL U1428 ( .A(b[10]), .B(n1004), .Y(n748) );
  XNOR2XL U1429 ( .A(b[12]), .B(n1006), .Y(n712) );
  XNOR2XL U1430 ( .A(b[11]), .B(n1004), .Y(n747) );
  XNOR2XL U1431 ( .A(b[15]), .B(n1006), .Y(n709) );
  XNOR2XL U1432 ( .A(b[13]), .B(n1005), .Y(n728) );
  XNOR2XL U1433 ( .A(b[14]), .B(n1006), .Y(n710) );
  NOR2X4 U1434 ( .A(n378), .B(n371), .Y(n183) );
  OAI22XL U1435 ( .A0(n24), .A1(n763), .B0(n762), .B1(n22), .Y(n630) );
  NOR2X4 U1436 ( .A(n389), .B(n398), .Y(n199) );
  INVX4 U1437 ( .A(n235), .Y(n234) );
  NAND2X2 U1438 ( .A(n209), .B(n221), .Y(n207) );
  NOR2X4 U1439 ( .A(n379), .B(n388), .Y(n188) );
  AOI21X4 U1440 ( .A0(n255), .A1(n236), .B0(n237), .Y(n235) );
  NOR2BXL U1441 ( .AN(b[0]), .B(n867), .Y(product[0]) );
  NOR2BXL U1442 ( .AN(b[0]), .B(n46), .Y(n579) );
  NOR2BXL U1443 ( .AN(b[0]), .B(n22), .Y(n643) );
  NOR2BXL U1444 ( .AN(b[0]), .B(n958), .Y(n627) );
  XNOR2X1 U1445 ( .A(b[0]), .B(n1001), .Y(n809) );
  NOR2BXL U1446 ( .AN(b[0]), .B(n34), .Y(n611) );
  NAND2BX1 U1447 ( .AN(b[0]), .B(n1004), .Y(n759) );
  NOR2BXL U1448 ( .AN(b[0]), .B(n961), .Y(n595) );
  NOR2BX1 U1449 ( .AN(b[0]), .B(n9), .Y(n675) );
  XNOR2X1 U1450 ( .A(b[0]), .B(n1005), .Y(n741) );
endmodule


module compare_1 ( clk, rst, sum, length );
  input [39:0] sum;
  output [5:0] length;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139;

  NAND2X1 U3 ( .A(n14), .B(n15), .Y(n110) );
  OAI2BB1X1 U4 ( .A0N(n3), .A1N(n137), .B0(n138), .Y(n125) );
  INVX2 U5 ( .A(n123), .Y(n3) );
  AOI31X1 U6 ( .A0(n122), .A1(n9), .A2(n121), .B0(n130), .Y(n123) );
  NAND4X1 U7 ( .A(n4), .B(n5), .C(n6), .D(n7), .Y(n122) );
  NAND4X1 U8 ( .A(n10), .B(n11), .C(n12), .D(n13), .Y(n130) );
  NAND4X1 U9 ( .A(n24), .B(n25), .C(n26), .D(n27), .Y(n131) );
  INVX2 U10 ( .A(n139), .Y(n21) );
  AOI31X1 U11 ( .A0(n139), .A1(n138), .A2(n137), .B0(length[5]), .Y(length[4])
         );
  NAND3X1 U12 ( .A(n30), .B(n31), .C(n127), .Y(n136) );
  OAI21X1 U13 ( .A0(n96), .A1(sum[24]), .B0(n22), .Y(n97) );
  AOI21X1 U14 ( .A0(n19), .A1(n95), .B0(sum[23]), .Y(n96) );
  OAI21X1 U15 ( .A0(n94), .A1(sum[20]), .B0(n18), .Y(n95) );
  AOI21X1 U16 ( .A0(n15), .A1(n93), .B0(sum[19]), .Y(n94) );
  OAI21X1 U17 ( .A0(n92), .A1(sum[16]), .B0(n14), .Y(n93) );
  AOI21X1 U18 ( .A0(n13), .A1(n91), .B0(sum[15]), .Y(n92) );
  OAI21X1 U19 ( .A0(n90), .A1(sum[12]), .B0(n12), .Y(n91) );
  AOI21X1 U20 ( .A0(n9), .A1(n89), .B0(sum[11]), .Y(n90) );
  OAI21X1 U21 ( .A0(n100), .A1(sum[32]), .B0(n28), .Y(n101) );
  AOI21X1 U22 ( .A0(n27), .A1(n99), .B0(sum[31]), .Y(n100) );
  OAI21X1 U23 ( .A0(n98), .A1(sum[28]), .B0(n26), .Y(n99) );
  AOI21X1 U24 ( .A0(n23), .A1(n97), .B0(sum[27]), .Y(n98) );
  OAI21X1 U25 ( .A0(n88), .A1(sum[8]), .B0(n8), .Y(n89) );
  AOI21X1 U26 ( .A0(n7), .A1(n87), .B0(sum[7]), .Y(n88) );
  OAI21X1 U27 ( .A0(n86), .A1(sum[4]), .B0(n6), .Y(n87) );
  AOI2BB1X1 U28 ( .A0N(n2), .A1N(sum[2]), .B0(sum[3]), .Y(n86) );
  AOI2BB1X1 U29 ( .A0N(sum[38]), .A1N(n103), .B0(sum[39]), .Y(length[0]) );
  AOI2BB1X1 U30 ( .A0N(n102), .A1N(sum[36]), .B0(sum[37]), .Y(n103) );
  AOI21X1 U31 ( .A0(n29), .A1(n101), .B0(sum[35]), .Y(n102) );
  INVX2 U32 ( .A(sum[1]), .Y(n2) );
  INVX2 U33 ( .A(sum[6]), .Y(n7) );
  AOI31X1 U34 ( .A0(n12), .A1(n13), .A2(n109), .B0(n108), .Y(n111) );
  OR2X1 U35 ( .A(sum[15]), .B(sum[16]), .Y(n108) );
  OAI211X1 U36 ( .A0(n107), .A1(n106), .B0(n10), .C0(n11), .Y(n109) );
  NAND2X1 U37 ( .A(n9), .B(n8), .Y(n106) );
  AOI31X1 U38 ( .A0(n18), .A1(n19), .A2(n113), .B0(n112), .Y(n115) );
  OR2X1 U39 ( .A(sum[23]), .B(sum[24]), .Y(n112) );
  OAI211X1 U40 ( .A0(n111), .A1(n110), .B0(n16), .C0(n17), .Y(n113) );
  INVX2 U41 ( .A(sum[20]), .Y(n17) );
  INVX2 U42 ( .A(sum[3]), .Y(n4) );
  AOI21X1 U43 ( .A0(n127), .A1(n120), .B0(sum[39]), .Y(length[1]) );
  OAI211X1 U44 ( .A0(n119), .A1(n118), .B0(n30), .C0(n31), .Y(n120) );
  NAND2X1 U45 ( .A(n28), .B(n29), .Y(n118) );
  AOI31X1 U46 ( .A0(n6), .A1(n7), .A2(n105), .B0(n104), .Y(n107) );
  OR2X1 U47 ( .A(sum[7]), .B(sum[8]), .Y(n104) );
  OAI211X1 U48 ( .A0(sum[1]), .A1(sum[2]), .B0(n4), .C0(n5), .Y(n105) );
  AOI31X1 U49 ( .A0(n26), .A1(n27), .A2(n117), .B0(n116), .Y(n119) );
  OR2X1 U50 ( .A(sum[31]), .B(sum[32]), .Y(n116) );
  OAI211X1 U51 ( .A0(n115), .A1(n114), .B0(n24), .C0(n25), .Y(n117) );
  NAND2X1 U52 ( .A(n22), .B(n23), .Y(n114) );
  INVX2 U53 ( .A(sum[4]), .Y(n5) );
  INVX2 U54 ( .A(sum[5]), .Y(n6) );
  INVX2 U55 ( .A(sum[10]), .Y(n9) );
  INVX2 U56 ( .A(sum[9]), .Y(n8) );
  INVX2 U57 ( .A(sum[11]), .Y(n10) );
  INVX2 U58 ( .A(sum[14]), .Y(n13) );
  INVX2 U59 ( .A(sum[12]), .Y(n11) );
  INVX2 U60 ( .A(sum[13]), .Y(n12) );
  INVX2 U61 ( .A(sum[18]), .Y(n15) );
  INVX2 U62 ( .A(sum[17]), .Y(n14) );
  INVX2 U63 ( .A(sum[19]), .Y(n16) );
  NOR3X1 U64 ( .A(sum[7]), .B(sum[9]), .C(sum[8]), .Y(n121) );
  AOI2BB1X1 U65 ( .A0N(n128), .A1N(n136), .B0(sum[39]), .Y(length[2]) );
  NOR2X1 U66 ( .A(n126), .B(n135), .Y(n128) );
  AOI31X1 U67 ( .A0(n125), .A1(n20), .A2(n124), .B0(n131), .Y(n126) );
  INVX2 U68 ( .A(sum[22]), .Y(n19) );
  INVX2 U69 ( .A(sum[21]), .Y(n18) );
  NAND4BBX1 U70 ( .AN(n130), .BN(sum[7]), .C(n9), .D(n129), .Y(n133) );
  NOR2X1 U71 ( .A(sum[9]), .B(sum[8]), .Y(n129) );
  OAI31X1 U72 ( .A0(n135), .A1(n134), .A2(n136), .B0(n1), .Y(length[3]) );
  INVX2 U73 ( .A(sum[39]), .Y(n1) );
  AOI31X1 U74 ( .A0(n138), .A1(n133), .A2(n137), .B0(n21), .Y(n134) );
  NOR4BX1 U75 ( .AN(n132), .B(n131), .C(sum[23]), .D(sum[24]), .Y(n139) );
  NOR2X1 U76 ( .A(sum[26]), .B(sum[25]), .Y(n132) );
  INVX2 U77 ( .A(sum[30]), .Y(n27) );
  INVX2 U78 ( .A(sum[26]), .Y(n23) );
  INVX2 U79 ( .A(sum[27]), .Y(n24) );
  INVX2 U80 ( .A(sum[25]), .Y(n22) );
  NOR4X1 U81 ( .A(sum[19]), .B(sum[20]), .C(sum[21]), .D(sum[22]), .Y(n138) );
  OR4X2 U82 ( .A(sum[31]), .B(sum[32]), .C(sum[33]), .D(sum[34]), .Y(n135) );
  OR3X2 U83 ( .A(n136), .B(sum[39]), .C(n135), .Y(length[5]) );
  NOR4X1 U84 ( .A(sum[15]), .B(sum[16]), .C(sum[17]), .D(sum[18]), .Y(n137) );
  INVX2 U85 ( .A(sum[28]), .Y(n25) );
  INVX2 U86 ( .A(sum[29]), .Y(n26) );
  NOR3X1 U87 ( .A(sum[24]), .B(sum[26]), .C(sum[25]), .Y(n124) );
  INVX2 U88 ( .A(sum[23]), .Y(n20) );
  NOR2X1 U89 ( .A(sum[38]), .B(sum[37]), .Y(n127) );
  INVX2 U90 ( .A(sum[35]), .Y(n30) );
  INVX2 U91 ( .A(sum[34]), .Y(n29) );
  INVX2 U92 ( .A(sum[33]), .Y(n28) );
  INVX2 U93 ( .A(sum[36]), .Y(n31) );
endmodule


module compare_2 ( clk, rst, sum, length );
  input [39:0] sum;
  output [5:0] length;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139;

  NAND2X1 U3 ( .A(n14), .B(n15), .Y(n110) );
  OAI2BB1X1 U4 ( .A0N(n3), .A1N(n137), .B0(n138), .Y(n125) );
  INVX2 U5 ( .A(n123), .Y(n3) );
  AOI31X1 U6 ( .A0(n122), .A1(n9), .A2(n121), .B0(n130), .Y(n123) );
  NAND4X1 U7 ( .A(n4), .B(n5), .C(n6), .D(n7), .Y(n122) );
  NAND4X1 U8 ( .A(n10), .B(n11), .C(n12), .D(n13), .Y(n130) );
  NAND4X1 U9 ( .A(n24), .B(n25), .C(n26), .D(n27), .Y(n131) );
  INVX2 U10 ( .A(n139), .Y(n21) );
  AOI31X1 U11 ( .A0(n139), .A1(n138), .A2(n137), .B0(length[5]), .Y(length[4])
         );
  NAND3X1 U12 ( .A(n30), .B(n31), .C(n127), .Y(n136) );
  OAI21X1 U13 ( .A0(n96), .A1(sum[24]), .B0(n22), .Y(n97) );
  AOI21X1 U14 ( .A0(n19), .A1(n95), .B0(sum[23]), .Y(n96) );
  OAI21X1 U15 ( .A0(n94), .A1(sum[20]), .B0(n18), .Y(n95) );
  AOI21X1 U16 ( .A0(n15), .A1(n93), .B0(sum[19]), .Y(n94) );
  OAI21X1 U17 ( .A0(n88), .A1(sum[8]), .B0(n8), .Y(n89) );
  AOI21X1 U18 ( .A0(n7), .A1(n87), .B0(sum[7]), .Y(n88) );
  OAI21X1 U19 ( .A0(n86), .A1(sum[4]), .B0(n6), .Y(n87) );
  AOI2BB1X1 U20 ( .A0N(n2), .A1N(sum[2]), .B0(sum[3]), .Y(n86) );
  OAI21X1 U21 ( .A0(n92), .A1(sum[16]), .B0(n14), .Y(n93) );
  AOI21X1 U22 ( .A0(n13), .A1(n91), .B0(sum[15]), .Y(n92) );
  OAI21X1 U23 ( .A0(n90), .A1(sum[12]), .B0(n12), .Y(n91) );
  AOI21X1 U24 ( .A0(n9), .A1(n89), .B0(sum[11]), .Y(n90) );
  OAI21X1 U25 ( .A0(n100), .A1(sum[32]), .B0(n28), .Y(n101) );
  AOI21X1 U26 ( .A0(n27), .A1(n99), .B0(sum[31]), .Y(n100) );
  OAI21X1 U27 ( .A0(n98), .A1(sum[28]), .B0(n26), .Y(n99) );
  AOI21X1 U28 ( .A0(n23), .A1(n97), .B0(sum[27]), .Y(n98) );
  AOI2BB1X1 U29 ( .A0N(sum[38]), .A1N(n103), .B0(sum[39]), .Y(length[0]) );
  AOI2BB1X1 U30 ( .A0N(n102), .A1N(sum[36]), .B0(sum[37]), .Y(n103) );
  AOI21X1 U31 ( .A0(n29), .A1(n101), .B0(sum[35]), .Y(n102) );
  INVX2 U32 ( .A(sum[1]), .Y(n2) );
  INVX2 U33 ( .A(sum[6]), .Y(n7) );
  AOI31X1 U34 ( .A0(n12), .A1(n13), .A2(n109), .B0(n108), .Y(n111) );
  OR2X1 U35 ( .A(sum[15]), .B(sum[16]), .Y(n108) );
  OAI211X1 U36 ( .A0(n107), .A1(n106), .B0(n10), .C0(n11), .Y(n109) );
  NAND2X1 U37 ( .A(n9), .B(n8), .Y(n106) );
  AOI31X1 U38 ( .A0(n18), .A1(n19), .A2(n113), .B0(n112), .Y(n115) );
  OR2X1 U39 ( .A(sum[23]), .B(sum[24]), .Y(n112) );
  OAI211X1 U40 ( .A0(n111), .A1(n110), .B0(n16), .C0(n17), .Y(n113) );
  INVX2 U41 ( .A(sum[20]), .Y(n17) );
  INVX2 U42 ( .A(sum[3]), .Y(n4) );
  AOI21X1 U43 ( .A0(n127), .A1(n120), .B0(sum[39]), .Y(length[1]) );
  OAI211X1 U44 ( .A0(n119), .A1(n118), .B0(n30), .C0(n31), .Y(n120) );
  NAND2X1 U45 ( .A(n28), .B(n29), .Y(n118) );
  AOI31X1 U46 ( .A0(n6), .A1(n7), .A2(n105), .B0(n104), .Y(n107) );
  OR2X1 U47 ( .A(sum[7]), .B(sum[8]), .Y(n104) );
  OAI211X1 U48 ( .A0(sum[1]), .A1(sum[2]), .B0(n4), .C0(n5), .Y(n105) );
  AOI31X1 U49 ( .A0(n26), .A1(n27), .A2(n117), .B0(n116), .Y(n119) );
  OR2X1 U50 ( .A(sum[31]), .B(sum[32]), .Y(n116) );
  OAI211X1 U51 ( .A0(n115), .A1(n114), .B0(n24), .C0(n25), .Y(n117) );
  NAND2X1 U52 ( .A(n22), .B(n23), .Y(n114) );
  INVX2 U53 ( .A(sum[5]), .Y(n6) );
  INVX2 U54 ( .A(sum[10]), .Y(n9) );
  INVX2 U55 ( .A(sum[4]), .Y(n5) );
  INVX2 U56 ( .A(sum[9]), .Y(n8) );
  INVX2 U57 ( .A(sum[14]), .Y(n13) );
  INVX2 U58 ( .A(sum[11]), .Y(n10) );
  INVX2 U59 ( .A(sum[13]), .Y(n12) );
  INVX2 U60 ( .A(sum[12]), .Y(n11) );
  INVX2 U61 ( .A(sum[18]), .Y(n15) );
  INVX2 U62 ( .A(sum[17]), .Y(n14) );
  NOR3X1 U63 ( .A(sum[7]), .B(sum[9]), .C(sum[8]), .Y(n121) );
  AOI2BB1X1 U64 ( .A0N(n128), .A1N(n136), .B0(sum[39]), .Y(length[2]) );
  NOR2X1 U65 ( .A(n126), .B(n135), .Y(n128) );
  AOI31X1 U66 ( .A0(n125), .A1(n20), .A2(n124), .B0(n131), .Y(n126) );
  INVX2 U67 ( .A(sum[22]), .Y(n19) );
  INVX2 U68 ( .A(sum[19]), .Y(n16) );
  INVX2 U69 ( .A(sum[21]), .Y(n18) );
  NAND4BBX1 U70 ( .AN(n130), .BN(sum[7]), .C(n9), .D(n129), .Y(n133) );
  NOR2X1 U71 ( .A(sum[9]), .B(sum[8]), .Y(n129) );
  OAI31X1 U72 ( .A0(n135), .A1(n134), .A2(n136), .B0(n1), .Y(length[3]) );
  INVX2 U73 ( .A(sum[39]), .Y(n1) );
  AOI31X1 U74 ( .A0(n138), .A1(n133), .A2(n137), .B0(n21), .Y(n134) );
  INVX2 U75 ( .A(sum[26]), .Y(n23) );
  INVX2 U76 ( .A(sum[25]), .Y(n22) );
  NOR4BX1 U77 ( .AN(n132), .B(n131), .C(sum[23]), .D(sum[24]), .Y(n139) );
  NOR2X1 U78 ( .A(sum[26]), .B(sum[25]), .Y(n132) );
  INVX2 U79 ( .A(sum[30]), .Y(n27) );
  INVX2 U80 ( .A(sum[27]), .Y(n24) );
  NOR4X1 U81 ( .A(sum[19]), .B(sum[20]), .C(sum[21]), .D(sum[22]), .Y(n138) );
  OR4X2 U82 ( .A(sum[31]), .B(sum[32]), .C(sum[33]), .D(sum[34]), .Y(n135) );
  OR3X2 U83 ( .A(n136), .B(sum[39]), .C(n135), .Y(length[5]) );
  NOR4X1 U84 ( .A(sum[15]), .B(sum[16]), .C(sum[17]), .D(sum[18]), .Y(n137) );
  INVX2 U85 ( .A(sum[28]), .Y(n25) );
  INVX2 U86 ( .A(sum[29]), .Y(n26) );
  NOR3X1 U87 ( .A(sum[24]), .B(sum[26]), .C(sum[25]), .Y(n124) );
  INVX2 U88 ( .A(sum[23]), .Y(n20) );
  NOR2X1 U89 ( .A(sum[38]), .B(sum[37]), .Y(n127) );
  INVX2 U90 ( .A(sum[35]), .Y(n30) );
  INVX2 U91 ( .A(sum[33]), .Y(n28) );
  INVX2 U92 ( .A(sum[34]), .Y(n29) );
  INVX2 U93 ( .A(sum[36]), .Y(n31) );
endmodule


module compare_3 ( clk, rst, sum, length );
  input [39:0] sum;
  output [5:0] length;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139;

  NAND2X1 U3 ( .A(n14), .B(n15), .Y(n110) );
  OAI2BB1X1 U4 ( .A0N(n3), .A1N(n137), .B0(n138), .Y(n125) );
  INVX2 U5 ( .A(n123), .Y(n3) );
  AOI31X1 U6 ( .A0(n122), .A1(n9), .A2(n121), .B0(n130), .Y(n123) );
  NAND4X1 U7 ( .A(n4), .B(n5), .C(n6), .D(n7), .Y(n122) );
  NAND4X1 U8 ( .A(n10), .B(n11), .C(n12), .D(n13), .Y(n130) );
  NAND4X1 U9 ( .A(n24), .B(n25), .C(n26), .D(n27), .Y(n131) );
  INVX2 U10 ( .A(n139), .Y(n21) );
  AOI31X1 U11 ( .A0(n139), .A1(n138), .A2(n137), .B0(length[5]), .Y(length[4])
         );
  NAND3X1 U12 ( .A(n30), .B(n31), .C(n127), .Y(n136) );
  OAI21X1 U13 ( .A0(n96), .A1(sum[24]), .B0(n22), .Y(n97) );
  AOI21X1 U14 ( .A0(n19), .A1(n95), .B0(sum[23]), .Y(n96) );
  OAI21X1 U15 ( .A0(n94), .A1(sum[20]), .B0(n18), .Y(n95) );
  AOI21X1 U16 ( .A0(n15), .A1(n93), .B0(sum[19]), .Y(n94) );
  OAI21X1 U17 ( .A0(n88), .A1(sum[8]), .B0(n8), .Y(n89) );
  AOI21X1 U18 ( .A0(n7), .A1(n87), .B0(sum[7]), .Y(n88) );
  OAI21X1 U19 ( .A0(n86), .A1(sum[4]), .B0(n6), .Y(n87) );
  AOI2BB1X1 U20 ( .A0N(n2), .A1N(sum[2]), .B0(sum[3]), .Y(n86) );
  OAI21X1 U21 ( .A0(n92), .A1(sum[16]), .B0(n14), .Y(n93) );
  AOI21X1 U22 ( .A0(n13), .A1(n91), .B0(sum[15]), .Y(n92) );
  OAI21X1 U23 ( .A0(n90), .A1(sum[12]), .B0(n12), .Y(n91) );
  AOI21X1 U24 ( .A0(n9), .A1(n89), .B0(sum[11]), .Y(n90) );
  OAI21X1 U25 ( .A0(n100), .A1(sum[32]), .B0(n28), .Y(n101) );
  AOI21X1 U26 ( .A0(n27), .A1(n99), .B0(sum[31]), .Y(n100) );
  OAI21X1 U27 ( .A0(n98), .A1(sum[28]), .B0(n26), .Y(n99) );
  AOI21X1 U28 ( .A0(n23), .A1(n97), .B0(sum[27]), .Y(n98) );
  AOI2BB1X1 U29 ( .A0N(sum[38]), .A1N(n103), .B0(sum[39]), .Y(length[0]) );
  AOI2BB1X1 U30 ( .A0N(n102), .A1N(sum[36]), .B0(sum[37]), .Y(n103) );
  AOI21X1 U31 ( .A0(n29), .A1(n101), .B0(sum[35]), .Y(n102) );
  INVX2 U32 ( .A(sum[1]), .Y(n2) );
  INVX2 U33 ( .A(sum[6]), .Y(n7) );
  AOI31X1 U34 ( .A0(n12), .A1(n13), .A2(n109), .B0(n108), .Y(n111) );
  OR2X1 U35 ( .A(sum[15]), .B(sum[16]), .Y(n108) );
  OAI211X1 U36 ( .A0(n107), .A1(n106), .B0(n10), .C0(n11), .Y(n109) );
  NAND2X1 U37 ( .A(n9), .B(n8), .Y(n106) );
  AOI31X1 U38 ( .A0(n18), .A1(n19), .A2(n113), .B0(n112), .Y(n115) );
  OR2X1 U39 ( .A(sum[23]), .B(sum[24]), .Y(n112) );
  OAI211X1 U40 ( .A0(n111), .A1(n110), .B0(n16), .C0(n17), .Y(n113) );
  INVX2 U41 ( .A(sum[20]), .Y(n17) );
  INVX2 U42 ( .A(sum[3]), .Y(n4) );
  AOI21X1 U43 ( .A0(n127), .A1(n120), .B0(sum[39]), .Y(length[1]) );
  OAI211X1 U44 ( .A0(n119), .A1(n118), .B0(n30), .C0(n31), .Y(n120) );
  NAND2X1 U45 ( .A(n28), .B(n29), .Y(n118) );
  AOI31X1 U46 ( .A0(n6), .A1(n7), .A2(n105), .B0(n104), .Y(n107) );
  OR2X1 U47 ( .A(sum[7]), .B(sum[8]), .Y(n104) );
  OAI211X1 U48 ( .A0(sum[1]), .A1(sum[2]), .B0(n4), .C0(n5), .Y(n105) );
  AOI31X1 U49 ( .A0(n26), .A1(n27), .A2(n117), .B0(n116), .Y(n119) );
  OR2X1 U50 ( .A(sum[31]), .B(sum[32]), .Y(n116) );
  OAI211X1 U51 ( .A0(n115), .A1(n114), .B0(n24), .C0(n25), .Y(n117) );
  NAND2X1 U52 ( .A(n22), .B(n23), .Y(n114) );
  INVX2 U53 ( .A(sum[5]), .Y(n6) );
  INVX2 U54 ( .A(sum[4]), .Y(n5) );
  INVX2 U55 ( .A(sum[10]), .Y(n9) );
  INVX2 U56 ( .A(sum[9]), .Y(n8) );
  INVX2 U57 ( .A(sum[11]), .Y(n10) );
  INVX2 U58 ( .A(sum[14]), .Y(n13) );
  INVX2 U59 ( .A(sum[13]), .Y(n12) );
  INVX2 U60 ( .A(sum[12]), .Y(n11) );
  INVX2 U61 ( .A(sum[18]), .Y(n15) );
  INVX2 U62 ( .A(sum[17]), .Y(n14) );
  INVX2 U63 ( .A(sum[19]), .Y(n16) );
  NOR3X1 U64 ( .A(sum[7]), .B(sum[9]), .C(sum[8]), .Y(n121) );
  AOI2BB1X1 U65 ( .A0N(n128), .A1N(n136), .B0(sum[39]), .Y(length[2]) );
  NOR2X1 U66 ( .A(n126), .B(n135), .Y(n128) );
  AOI31X1 U67 ( .A0(n125), .A1(n20), .A2(n124), .B0(n131), .Y(n126) );
  INVX2 U68 ( .A(sum[22]), .Y(n19) );
  INVX2 U69 ( .A(sum[21]), .Y(n18) );
  NAND4BBX1 U70 ( .AN(n130), .BN(sum[7]), .C(n9), .D(n129), .Y(n133) );
  NOR2X1 U71 ( .A(sum[9]), .B(sum[8]), .Y(n129) );
  OAI31X1 U72 ( .A0(n135), .A1(n134), .A2(n136), .B0(n1), .Y(length[3]) );
  INVX2 U73 ( .A(sum[39]), .Y(n1) );
  AOI31X1 U74 ( .A0(n138), .A1(n133), .A2(n137), .B0(n21), .Y(n134) );
  INVX2 U75 ( .A(sum[26]), .Y(n23) );
  INVX2 U76 ( .A(sum[25]), .Y(n22) );
  NOR4BX1 U77 ( .AN(n132), .B(n131), .C(sum[23]), .D(sum[24]), .Y(n139) );
  NOR2X1 U78 ( .A(sum[26]), .B(sum[25]), .Y(n132) );
  INVX2 U79 ( .A(sum[30]), .Y(n27) );
  INVX2 U80 ( .A(sum[27]), .Y(n24) );
  NOR4X1 U81 ( .A(sum[19]), .B(sum[20]), .C(sum[21]), .D(sum[22]), .Y(n138) );
  OR4X2 U82 ( .A(sum[31]), .B(sum[32]), .C(sum[33]), .D(sum[34]), .Y(n135) );
  OR3X2 U83 ( .A(n136), .B(sum[39]), .C(n135), .Y(length[5]) );
  NOR4X1 U84 ( .A(sum[15]), .B(sum[16]), .C(sum[17]), .D(sum[18]), .Y(n137) );
  INVX2 U85 ( .A(sum[28]), .Y(n25) );
  INVX2 U86 ( .A(sum[29]), .Y(n26) );
  NOR3X1 U87 ( .A(sum[24]), .B(sum[26]), .C(sum[25]), .Y(n124) );
  INVX2 U88 ( .A(sum[23]), .Y(n20) );
  NOR2X1 U89 ( .A(sum[38]), .B(sum[37]), .Y(n127) );
  INVX2 U90 ( .A(sum[35]), .Y(n30) );
  INVX2 U91 ( .A(sum[33]), .Y(n28) );
  INVX2 U92 ( .A(sum[34]), .Y(n29) );
  INVX2 U93 ( .A(sum[36]), .Y(n31) );
endmodule


module compare_4 ( clk, rst, sum, length );
  input [39:0] sum;
  output [5:0] length;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139;

  NAND2X1 U3 ( .A(n14), .B(n15), .Y(n110) );
  OAI2BB1X1 U4 ( .A0N(n3), .A1N(n137), .B0(n138), .Y(n125) );
  INVX2 U5 ( .A(n123), .Y(n3) );
  AOI31X1 U6 ( .A0(n122), .A1(n9), .A2(n121), .B0(n130), .Y(n123) );
  NAND4X1 U7 ( .A(n4), .B(n5), .C(n6), .D(n7), .Y(n122) );
  NAND4X1 U8 ( .A(n10), .B(n11), .C(n12), .D(n13), .Y(n130) );
  NAND4X1 U9 ( .A(n24), .B(n25), .C(n26), .D(n27), .Y(n131) );
  INVX2 U10 ( .A(n139), .Y(n21) );
  AOI31X1 U11 ( .A0(n139), .A1(n138), .A2(n137), .B0(length[5]), .Y(length[4])
         );
  NAND3X1 U12 ( .A(n30), .B(n31), .C(n127), .Y(n136) );
  OAI21X1 U13 ( .A0(n96), .A1(sum[24]), .B0(n22), .Y(n97) );
  AOI21X1 U14 ( .A0(n19), .A1(n95), .B0(sum[23]), .Y(n96) );
  OAI21X1 U15 ( .A0(n94), .A1(sum[20]), .B0(n18), .Y(n95) );
  AOI21X1 U16 ( .A0(n15), .A1(n93), .B0(sum[19]), .Y(n94) );
  OAI21X1 U17 ( .A0(n88), .A1(sum[8]), .B0(n8), .Y(n89) );
  AOI21X1 U18 ( .A0(n7), .A1(n87), .B0(sum[7]), .Y(n88) );
  OAI21X1 U19 ( .A0(n86), .A1(sum[4]), .B0(n6), .Y(n87) );
  AOI2BB1X1 U20 ( .A0N(n2), .A1N(sum[2]), .B0(sum[3]), .Y(n86) );
  OAI21X1 U21 ( .A0(n92), .A1(sum[16]), .B0(n14), .Y(n93) );
  AOI21X1 U22 ( .A0(n13), .A1(n91), .B0(sum[15]), .Y(n92) );
  OAI21X1 U23 ( .A0(n90), .A1(sum[12]), .B0(n12), .Y(n91) );
  AOI21X1 U24 ( .A0(n9), .A1(n89), .B0(sum[11]), .Y(n90) );
  OAI21X1 U25 ( .A0(n100), .A1(sum[32]), .B0(n28), .Y(n101) );
  AOI21X1 U26 ( .A0(n27), .A1(n99), .B0(sum[31]), .Y(n100) );
  OAI21X1 U27 ( .A0(n98), .A1(sum[28]), .B0(n26), .Y(n99) );
  AOI21X1 U28 ( .A0(n23), .A1(n97), .B0(sum[27]), .Y(n98) );
  AOI2BB1X1 U29 ( .A0N(sum[38]), .A1N(n103), .B0(sum[39]), .Y(length[0]) );
  AOI2BB1X1 U30 ( .A0N(n102), .A1N(sum[36]), .B0(sum[37]), .Y(n103) );
  AOI21X1 U31 ( .A0(n29), .A1(n101), .B0(sum[35]), .Y(n102) );
  INVX2 U32 ( .A(sum[1]), .Y(n2) );
  INVX2 U33 ( .A(sum[6]), .Y(n7) );
  AOI31X1 U34 ( .A0(n12), .A1(n13), .A2(n109), .B0(n108), .Y(n111) );
  OR2X1 U35 ( .A(sum[15]), .B(sum[16]), .Y(n108) );
  OAI211X1 U36 ( .A0(n107), .A1(n106), .B0(n10), .C0(n11), .Y(n109) );
  NAND2X1 U37 ( .A(n9), .B(n8), .Y(n106) );
  AOI31X1 U38 ( .A0(n18), .A1(n19), .A2(n113), .B0(n112), .Y(n115) );
  OR2X1 U39 ( .A(sum[23]), .B(sum[24]), .Y(n112) );
  OAI211X1 U40 ( .A0(n111), .A1(n110), .B0(n16), .C0(n17), .Y(n113) );
  INVX2 U41 ( .A(sum[20]), .Y(n17) );
  INVX2 U42 ( .A(sum[3]), .Y(n4) );
  AOI21X1 U43 ( .A0(n127), .A1(n120), .B0(sum[39]), .Y(length[1]) );
  OAI211X1 U44 ( .A0(n119), .A1(n118), .B0(n30), .C0(n31), .Y(n120) );
  NAND2X1 U45 ( .A(n28), .B(n29), .Y(n118) );
  AOI31X1 U46 ( .A0(n6), .A1(n7), .A2(n105), .B0(n104), .Y(n107) );
  OR2X1 U47 ( .A(sum[7]), .B(sum[8]), .Y(n104) );
  OAI211X1 U48 ( .A0(sum[1]), .A1(sum[2]), .B0(n4), .C0(n5), .Y(n105) );
  AOI31X1 U49 ( .A0(n26), .A1(n27), .A2(n117), .B0(n116), .Y(n119) );
  OR2X1 U50 ( .A(sum[31]), .B(sum[32]), .Y(n116) );
  OAI211X1 U51 ( .A0(n115), .A1(n114), .B0(n24), .C0(n25), .Y(n117) );
  NAND2X1 U52 ( .A(n22), .B(n23), .Y(n114) );
  INVX2 U53 ( .A(sum[5]), .Y(n6) );
  INVX2 U54 ( .A(sum[4]), .Y(n5) );
  INVX2 U55 ( .A(sum[10]), .Y(n9) );
  INVX2 U56 ( .A(sum[9]), .Y(n8) );
  INVX2 U57 ( .A(sum[11]), .Y(n10) );
  INVX2 U58 ( .A(sum[14]), .Y(n13) );
  INVX2 U59 ( .A(sum[13]), .Y(n12) );
  INVX2 U60 ( .A(sum[12]), .Y(n11) );
  INVX2 U61 ( .A(sum[18]), .Y(n15) );
  INVX2 U62 ( .A(sum[17]), .Y(n14) );
  INVX2 U63 ( .A(sum[19]), .Y(n16) );
  NOR3X1 U64 ( .A(sum[7]), .B(sum[9]), .C(sum[8]), .Y(n121) );
  AOI2BB1X1 U65 ( .A0N(n128), .A1N(n136), .B0(sum[39]), .Y(length[2]) );
  NOR2X1 U66 ( .A(n126), .B(n135), .Y(n128) );
  AOI31X1 U67 ( .A0(n125), .A1(n20), .A2(n124), .B0(n131), .Y(n126) );
  INVX2 U68 ( .A(sum[22]), .Y(n19) );
  INVX2 U69 ( .A(sum[21]), .Y(n18) );
  NAND4BBX1 U70 ( .AN(n130), .BN(sum[7]), .C(n9), .D(n129), .Y(n133) );
  NOR2X1 U71 ( .A(sum[9]), .B(sum[8]), .Y(n129) );
  OAI31X1 U72 ( .A0(n135), .A1(n134), .A2(n136), .B0(n1), .Y(length[3]) );
  INVX2 U73 ( .A(sum[39]), .Y(n1) );
  AOI31X1 U74 ( .A0(n138), .A1(n133), .A2(n137), .B0(n21), .Y(n134) );
  INVX2 U75 ( .A(sum[26]), .Y(n23) );
  INVX2 U76 ( .A(sum[25]), .Y(n22) );
  NOR4BX1 U77 ( .AN(n132), .B(n131), .C(sum[23]), .D(sum[24]), .Y(n139) );
  NOR2X1 U78 ( .A(sum[26]), .B(sum[25]), .Y(n132) );
  INVX2 U79 ( .A(sum[30]), .Y(n27) );
  INVX2 U80 ( .A(sum[27]), .Y(n24) );
  NOR4X1 U81 ( .A(sum[19]), .B(sum[20]), .C(sum[21]), .D(sum[22]), .Y(n138) );
  OR4X2 U82 ( .A(sum[31]), .B(sum[32]), .C(sum[33]), .D(sum[34]), .Y(n135) );
  OR3X2 U83 ( .A(n136), .B(sum[39]), .C(n135), .Y(length[5]) );
  NOR4X1 U84 ( .A(sum[15]), .B(sum[16]), .C(sum[17]), .D(sum[18]), .Y(n137) );
  INVX2 U85 ( .A(sum[28]), .Y(n25) );
  INVX2 U86 ( .A(sum[29]), .Y(n26) );
  NOR3X1 U87 ( .A(sum[24]), .B(sum[26]), .C(sum[25]), .Y(n124) );
  INVX2 U88 ( .A(sum[23]), .Y(n20) );
  NOR2X1 U89 ( .A(sum[38]), .B(sum[37]), .Y(n127) );
  INVX2 U90 ( .A(sum[35]), .Y(n30) );
  INVX2 U91 ( .A(sum[33]), .Y(n28) );
  INVX2 U92 ( .A(sum[34]), .Y(n29) );
  INVX2 U93 ( .A(sum[36]), .Y(n31) );
endmodule


module compare_5 ( clk, rst, sum, length );
  input [39:0] sum;
  output [5:0] length;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139;

  NAND2X1 U3 ( .A(n14), .B(n15), .Y(n110) );
  OAI2BB1X1 U4 ( .A0N(n3), .A1N(n137), .B0(n138), .Y(n125) );
  INVX2 U5 ( .A(n123), .Y(n3) );
  AOI31X1 U6 ( .A0(n122), .A1(n9), .A2(n121), .B0(n130), .Y(n123) );
  NAND4X1 U7 ( .A(n4), .B(n5), .C(n6), .D(n7), .Y(n122) );
  NAND4X1 U8 ( .A(n10), .B(n11), .C(n12), .D(n13), .Y(n130) );
  NAND4X1 U9 ( .A(n24), .B(n25), .C(n26), .D(n27), .Y(n131) );
  INVX2 U10 ( .A(n139), .Y(n21) );
  AOI31X1 U11 ( .A0(n139), .A1(n138), .A2(n137), .B0(length[5]), .Y(length[4])
         );
  NAND3X1 U12 ( .A(n30), .B(n31), .C(n127), .Y(n136) );
  OAI21X1 U13 ( .A0(n96), .A1(sum[24]), .B0(n22), .Y(n97) );
  AOI21X1 U14 ( .A0(n19), .A1(n95), .B0(sum[23]), .Y(n96) );
  OAI21X1 U15 ( .A0(n94), .A1(sum[20]), .B0(n18), .Y(n95) );
  AOI21X1 U16 ( .A0(n15), .A1(n93), .B0(sum[19]), .Y(n94) );
  OAI21X1 U17 ( .A0(n88), .A1(sum[8]), .B0(n8), .Y(n89) );
  AOI21X1 U18 ( .A0(n7), .A1(n87), .B0(sum[7]), .Y(n88) );
  OAI21X1 U19 ( .A0(n86), .A1(sum[4]), .B0(n6), .Y(n87) );
  AOI2BB1X1 U20 ( .A0N(n2), .A1N(sum[2]), .B0(sum[3]), .Y(n86) );
  OAI21X1 U21 ( .A0(n92), .A1(sum[16]), .B0(n14), .Y(n93) );
  AOI21X1 U22 ( .A0(n13), .A1(n91), .B0(sum[15]), .Y(n92) );
  OAI21X1 U23 ( .A0(n90), .A1(sum[12]), .B0(n12), .Y(n91) );
  AOI21X1 U24 ( .A0(n9), .A1(n89), .B0(sum[11]), .Y(n90) );
  OAI21X1 U25 ( .A0(n100), .A1(sum[32]), .B0(n28), .Y(n101) );
  AOI21X1 U26 ( .A0(n27), .A1(n99), .B0(sum[31]), .Y(n100) );
  OAI21X1 U27 ( .A0(n98), .A1(sum[28]), .B0(n26), .Y(n99) );
  AOI21X1 U28 ( .A0(n23), .A1(n97), .B0(sum[27]), .Y(n98) );
  AOI2BB1X1 U29 ( .A0N(sum[38]), .A1N(n103), .B0(sum[39]), .Y(length[0]) );
  AOI2BB1X1 U30 ( .A0N(n102), .A1N(sum[36]), .B0(sum[37]), .Y(n103) );
  AOI21X1 U31 ( .A0(n29), .A1(n101), .B0(sum[35]), .Y(n102) );
  INVX2 U32 ( .A(sum[1]), .Y(n2) );
  INVX2 U33 ( .A(sum[6]), .Y(n7) );
  AOI31X1 U34 ( .A0(n12), .A1(n13), .A2(n109), .B0(n108), .Y(n111) );
  OR2X1 U35 ( .A(sum[15]), .B(sum[16]), .Y(n108) );
  OAI211X1 U36 ( .A0(n107), .A1(n106), .B0(n10), .C0(n11), .Y(n109) );
  NAND2X1 U37 ( .A(n9), .B(n8), .Y(n106) );
  AOI31X1 U38 ( .A0(n18), .A1(n19), .A2(n113), .B0(n112), .Y(n115) );
  OR2X1 U39 ( .A(sum[23]), .B(sum[24]), .Y(n112) );
  OAI211X1 U40 ( .A0(n111), .A1(n110), .B0(n16), .C0(n17), .Y(n113) );
  INVX2 U41 ( .A(sum[20]), .Y(n17) );
  INVX2 U42 ( .A(sum[3]), .Y(n4) );
  AOI21X1 U43 ( .A0(n127), .A1(n120), .B0(sum[39]), .Y(length[1]) );
  OAI211X1 U44 ( .A0(n119), .A1(n118), .B0(n30), .C0(n31), .Y(n120) );
  NAND2X1 U45 ( .A(n28), .B(n29), .Y(n118) );
  AOI31X1 U46 ( .A0(n6), .A1(n7), .A2(n105), .B0(n104), .Y(n107) );
  OR2X1 U47 ( .A(sum[7]), .B(sum[8]), .Y(n104) );
  OAI211X1 U48 ( .A0(sum[1]), .A1(sum[2]), .B0(n4), .C0(n5), .Y(n105) );
  AOI31X1 U49 ( .A0(n26), .A1(n27), .A2(n117), .B0(n116), .Y(n119) );
  OR2X1 U50 ( .A(sum[31]), .B(sum[32]), .Y(n116) );
  OAI211X1 U51 ( .A0(n115), .A1(n114), .B0(n24), .C0(n25), .Y(n117) );
  NAND2X1 U52 ( .A(n22), .B(n23), .Y(n114) );
  INVX2 U53 ( .A(sum[5]), .Y(n6) );
  INVX2 U54 ( .A(sum[4]), .Y(n5) );
  INVX2 U55 ( .A(sum[10]), .Y(n9) );
  INVX2 U56 ( .A(sum[9]), .Y(n8) );
  INVX2 U57 ( .A(sum[11]), .Y(n10) );
  INVX2 U58 ( .A(sum[14]), .Y(n13) );
  INVX2 U59 ( .A(sum[13]), .Y(n12) );
  INVX2 U60 ( .A(sum[12]), .Y(n11) );
  INVX2 U61 ( .A(sum[18]), .Y(n15) );
  INVX2 U62 ( .A(sum[17]), .Y(n14) );
  INVX2 U63 ( .A(sum[19]), .Y(n16) );
  AOI2BB1X1 U64 ( .A0N(n128), .A1N(n136), .B0(sum[39]), .Y(length[2]) );
  NOR2X1 U65 ( .A(n126), .B(n135), .Y(n128) );
  AOI31X1 U66 ( .A0(n125), .A1(n20), .A2(n124), .B0(n131), .Y(n126) );
  NOR3X1 U67 ( .A(sum[7]), .B(sum[9]), .C(sum[8]), .Y(n121) );
  INVX2 U68 ( .A(sum[22]), .Y(n19) );
  INVX2 U69 ( .A(sum[21]), .Y(n18) );
  NAND4BBX1 U70 ( .AN(n130), .BN(sum[7]), .C(n9), .D(n129), .Y(n133) );
  NOR2X1 U71 ( .A(sum[9]), .B(sum[8]), .Y(n129) );
  OAI31X1 U72 ( .A0(n135), .A1(n134), .A2(n136), .B0(n1), .Y(length[3]) );
  INVX2 U73 ( .A(sum[39]), .Y(n1) );
  AOI31X1 U74 ( .A0(n138), .A1(n133), .A2(n137), .B0(n21), .Y(n134) );
  INVX2 U75 ( .A(sum[26]), .Y(n23) );
  INVX2 U76 ( .A(sum[25]), .Y(n22) );
  NOR4BX1 U77 ( .AN(n132), .B(n131), .C(sum[23]), .D(sum[24]), .Y(n139) );
  NOR2X1 U78 ( .A(sum[26]), .B(sum[25]), .Y(n132) );
  INVX2 U79 ( .A(sum[30]), .Y(n27) );
  INVX2 U80 ( .A(sum[27]), .Y(n24) );
  OR4X2 U81 ( .A(sum[31]), .B(sum[32]), .C(sum[33]), .D(sum[34]), .Y(n135) );
  OR3X2 U82 ( .A(n136), .B(sum[39]), .C(n135), .Y(length[5]) );
  NOR4X1 U83 ( .A(sum[19]), .B(sum[20]), .C(sum[21]), .D(sum[22]), .Y(n138) );
  NOR4X1 U84 ( .A(sum[15]), .B(sum[16]), .C(sum[17]), .D(sum[18]), .Y(n137) );
  INVX2 U85 ( .A(sum[28]), .Y(n25) );
  INVX2 U86 ( .A(sum[29]), .Y(n26) );
  NOR3X1 U87 ( .A(sum[24]), .B(sum[26]), .C(sum[25]), .Y(n124) );
  INVX2 U88 ( .A(sum[23]), .Y(n20) );
  NOR2X1 U89 ( .A(sum[38]), .B(sum[37]), .Y(n127) );
  INVX2 U90 ( .A(sum[35]), .Y(n30) );
  INVX2 U91 ( .A(sum[33]), .Y(n28) );
  INVX2 U92 ( .A(sum[34]), .Y(n29) );
  INVX2 U93 ( .A(sum[36]), .Y(n31) );
endmodule


module compare_6 ( clk, rst, sum, length );
  input [39:0] sum;
  output [5:0] length;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139;

  NAND2X1 U3 ( .A(n14), .B(n15), .Y(n110) );
  OAI2BB1X1 U4 ( .A0N(n3), .A1N(n137), .B0(n138), .Y(n125) );
  INVX2 U5 ( .A(n123), .Y(n3) );
  AOI31X1 U6 ( .A0(n122), .A1(n9), .A2(n121), .B0(n130), .Y(n123) );
  NAND4X1 U7 ( .A(n4), .B(n5), .C(n6), .D(n7), .Y(n122) );
  NAND4X1 U8 ( .A(n10), .B(n11), .C(n12), .D(n13), .Y(n130) );
  AOI31X1 U9 ( .A0(n139), .A1(n138), .A2(n137), .B0(length[5]), .Y(length[4])
         );
  NAND4X1 U10 ( .A(n24), .B(n25), .C(n26), .D(n27), .Y(n131) );
  INVX2 U11 ( .A(n139), .Y(n21) );
  NAND3X1 U12 ( .A(n30), .B(n31), .C(n127), .Y(n136) );
  AOI2BB1X1 U13 ( .A0N(sum[38]), .A1N(n103), .B0(sum[39]), .Y(length[0]) );
  AOI2BB1X1 U14 ( .A0N(n102), .A1N(sum[36]), .B0(sum[37]), .Y(n103) );
  AOI21X1 U15 ( .A0(n29), .A1(n101), .B0(sum[35]), .Y(n102) );
  OAI21X1 U16 ( .A0(n96), .A1(sum[24]), .B0(n22), .Y(n97) );
  AOI21X1 U17 ( .A0(n19), .A1(n95), .B0(sum[23]), .Y(n96) );
  OAI21X1 U18 ( .A0(n94), .A1(sum[20]), .B0(n18), .Y(n95) );
  AOI21X1 U19 ( .A0(n15), .A1(n93), .B0(sum[19]), .Y(n94) );
  OAI21X1 U20 ( .A0(n88), .A1(sum[8]), .B0(n8), .Y(n89) );
  AOI21X1 U21 ( .A0(n7), .A1(n87), .B0(sum[7]), .Y(n88) );
  OAI21X1 U22 ( .A0(n86), .A1(sum[4]), .B0(n6), .Y(n87) );
  AOI2BB1X1 U23 ( .A0N(n2), .A1N(sum[2]), .B0(sum[3]), .Y(n86) );
  OAI21X1 U24 ( .A0(n100), .A1(sum[32]), .B0(n28), .Y(n101) );
  AOI21X1 U25 ( .A0(n27), .A1(n99), .B0(sum[31]), .Y(n100) );
  OAI21X1 U26 ( .A0(n98), .A1(sum[28]), .B0(n26), .Y(n99) );
  AOI21X1 U27 ( .A0(n23), .A1(n97), .B0(sum[27]), .Y(n98) );
  OAI21X1 U28 ( .A0(n92), .A1(sum[16]), .B0(n14), .Y(n93) );
  AOI21X1 U29 ( .A0(n13), .A1(n91), .B0(sum[15]), .Y(n92) );
  OAI21X1 U30 ( .A0(n90), .A1(sum[12]), .B0(n12), .Y(n91) );
  AOI21X1 U31 ( .A0(n9), .A1(n89), .B0(sum[11]), .Y(n90) );
  INVX2 U32 ( .A(sum[1]), .Y(n2) );
  OAI211X1 U33 ( .A0(n119), .A1(n118), .B0(n30), .C0(n31), .Y(n120) );
  NAND2X1 U34 ( .A(n28), .B(n29), .Y(n118) );
  AOI31X1 U35 ( .A0(n6), .A1(n7), .A2(n105), .B0(n104), .Y(n107) );
  OR2X1 U36 ( .A(sum[7]), .B(sum[8]), .Y(n104) );
  OAI211X1 U37 ( .A0(sum[1]), .A1(sum[2]), .B0(n4), .C0(n5), .Y(n105) );
  AOI31X1 U38 ( .A0(n12), .A1(n13), .A2(n109), .B0(n108), .Y(n111) );
  OR2X1 U39 ( .A(sum[15]), .B(sum[16]), .Y(n108) );
  OAI211X1 U40 ( .A0(n107), .A1(n106), .B0(n10), .C0(n11), .Y(n109) );
  NAND2X1 U41 ( .A(n9), .B(n8), .Y(n106) );
  AOI31X1 U42 ( .A0(n18), .A1(n19), .A2(n113), .B0(n112), .Y(n115) );
  OR2X1 U43 ( .A(sum[23]), .B(sum[24]), .Y(n112) );
  OAI211X1 U44 ( .A0(n111), .A1(n110), .B0(n16), .C0(n17), .Y(n113) );
  INVX2 U45 ( .A(sum[20]), .Y(n17) );
  AOI31X1 U46 ( .A0(n26), .A1(n27), .A2(n117), .B0(n116), .Y(n119) );
  OR2X1 U47 ( .A(sum[31]), .B(sum[32]), .Y(n116) );
  OAI211X1 U48 ( .A0(n115), .A1(n114), .B0(n24), .C0(n25), .Y(n117) );
  NAND2X1 U49 ( .A(n22), .B(n23), .Y(n114) );
  INVX2 U50 ( .A(sum[3]), .Y(n4) );
  INVX2 U51 ( .A(sum[6]), .Y(n7) );
  INVX2 U52 ( .A(sum[5]), .Y(n6) );
  INVX2 U53 ( .A(sum[4]), .Y(n5) );
  INVX2 U54 ( .A(sum[10]), .Y(n9) );
  INVX2 U55 ( .A(sum[9]), .Y(n8) );
  INVX2 U56 ( .A(sum[11]), .Y(n10) );
  INVX2 U57 ( .A(sum[14]), .Y(n13) );
  INVX2 U58 ( .A(sum[13]), .Y(n12) );
  INVX2 U59 ( .A(sum[12]), .Y(n11) );
  INVX2 U60 ( .A(sum[18]), .Y(n15) );
  INVX2 U61 ( .A(sum[17]), .Y(n14) );
  INVX2 U62 ( .A(sum[19]), .Y(n16) );
  INVX2 U63 ( .A(sum[22]), .Y(n19) );
  NOR3X1 U64 ( .A(sum[7]), .B(sum[9]), .C(sum[8]), .Y(n121) );
  AOI2BB1X1 U65 ( .A0N(n128), .A1N(n136), .B0(sum[39]), .Y(length[2]) );
  NOR2X1 U66 ( .A(n126), .B(n135), .Y(n128) );
  AOI31X1 U67 ( .A0(n125), .A1(n20), .A2(n124), .B0(n131), .Y(n126) );
  INVX2 U68 ( .A(sum[21]), .Y(n18) );
  INVX2 U69 ( .A(sum[26]), .Y(n23) );
  NAND4BBX1 U70 ( .AN(n130), .BN(sum[7]), .C(n9), .D(n129), .Y(n133) );
  NOR2X1 U71 ( .A(sum[9]), .B(sum[8]), .Y(n129) );
  OAI31X1 U72 ( .A0(n135), .A1(n134), .A2(n136), .B0(n1), .Y(length[3]) );
  AOI31X1 U73 ( .A0(n138), .A1(n133), .A2(n137), .B0(n21), .Y(n134) );
  INVX2 U74 ( .A(sum[25]), .Y(n22) );
  NOR4BX1 U75 ( .AN(n132), .B(n131), .C(sum[23]), .D(sum[24]), .Y(n139) );
  NOR2X1 U76 ( .A(sum[26]), .B(sum[25]), .Y(n132) );
  INVX2 U77 ( .A(sum[30]), .Y(n27) );
  INVX2 U78 ( .A(sum[27]), .Y(n24) );
  OR4X2 U79 ( .A(sum[31]), .B(sum[32]), .C(sum[33]), .D(sum[34]), .Y(n135) );
  NOR4X1 U80 ( .A(sum[15]), .B(sum[16]), .C(sum[17]), .D(sum[18]), .Y(n137) );
  NOR4X1 U81 ( .A(sum[19]), .B(sum[20]), .C(sum[21]), .D(sum[22]), .Y(n138) );
  NOR3X1 U82 ( .A(sum[24]), .B(sum[26]), .C(sum[25]), .Y(n124) );
  INVX2 U83 ( .A(sum[28]), .Y(n25) );
  INVX2 U84 ( .A(sum[29]), .Y(n26) );
  INVX2 U85 ( .A(sum[23]), .Y(n20) );
  NOR2X1 U86 ( .A(sum[38]), .B(sum[37]), .Y(n127) );
  INVX2 U87 ( .A(sum[35]), .Y(n30) );
  INVX2 U88 ( .A(sum[34]), .Y(n29) );
  INVX2 U89 ( .A(sum[33]), .Y(n28) );
  INVX2 U90 ( .A(sum[36]), .Y(n31) );
  OR3X2 U91 ( .A(n136), .B(sum[39]), .C(n135), .Y(length[5]) );
  INVX2 U92 ( .A(sum[39]), .Y(n1) );
  AOI21X1 U93 ( .A0(n127), .A1(n120), .B0(sum[39]), .Y(length[1]) );
endmodule


module compare_7 ( clk, rst, sum, length );
  input [39:0] sum;
  output [5:0] length;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139;

  NAND2X1 U3 ( .A(n14), .B(n15), .Y(n110) );
  OAI2BB1X1 U4 ( .A0N(n3), .A1N(n137), .B0(n138), .Y(n125) );
  INVX2 U5 ( .A(n123), .Y(n3) );
  AOI31X1 U6 ( .A0(n122), .A1(n9), .A2(n121), .B0(n130), .Y(n123) );
  NAND4X1 U7 ( .A(n4), .B(n5), .C(n6), .D(n7), .Y(n122) );
  NAND4X1 U8 ( .A(n10), .B(n11), .C(n12), .D(n13), .Y(n130) );
  NAND4X1 U9 ( .A(n24), .B(n25), .C(n26), .D(n27), .Y(n131) );
  INVX2 U10 ( .A(n139), .Y(n21) );
  AOI31X1 U11 ( .A0(n139), .A1(n138), .A2(n137), .B0(length[5]), .Y(length[4])
         );
  NAND3X1 U12 ( .A(n30), .B(n31), .C(n127), .Y(n136) );
  OAI21X1 U13 ( .A0(n96), .A1(sum[24]), .B0(n22), .Y(n97) );
  AOI21X1 U14 ( .A0(n19), .A1(n95), .B0(sum[23]), .Y(n96) );
  OAI21X1 U15 ( .A0(n94), .A1(sum[20]), .B0(n18), .Y(n95) );
  AOI21X1 U16 ( .A0(n15), .A1(n93), .B0(sum[19]), .Y(n94) );
  OAI21X1 U17 ( .A0(n100), .A1(sum[32]), .B0(n28), .Y(n101) );
  AOI21X1 U18 ( .A0(n27), .A1(n99), .B0(sum[31]), .Y(n100) );
  OAI21X1 U19 ( .A0(n98), .A1(sum[28]), .B0(n26), .Y(n99) );
  AOI21X1 U20 ( .A0(n23), .A1(n97), .B0(sum[27]), .Y(n98) );
  OAI21X1 U21 ( .A0(n92), .A1(sum[16]), .B0(n14), .Y(n93) );
  AOI21X1 U22 ( .A0(n13), .A1(n91), .B0(sum[15]), .Y(n92) );
  OAI21X1 U23 ( .A0(n90), .A1(sum[12]), .B0(n12), .Y(n91) );
  AOI21X1 U24 ( .A0(n9), .A1(n89), .B0(sum[11]), .Y(n90) );
  OAI21X1 U25 ( .A0(n88), .A1(sum[8]), .B0(n8), .Y(n89) );
  AOI21X1 U26 ( .A0(n7), .A1(n87), .B0(sum[7]), .Y(n88) );
  OAI21X1 U27 ( .A0(n86), .A1(sum[4]), .B0(n6), .Y(n87) );
  AOI2BB1X1 U28 ( .A0N(n2), .A1N(sum[2]), .B0(sum[3]), .Y(n86) );
  AOI2BB1X1 U29 ( .A0N(sum[38]), .A1N(n103), .B0(sum[39]), .Y(length[0]) );
  AOI2BB1X1 U30 ( .A0N(n102), .A1N(sum[36]), .B0(sum[37]), .Y(n103) );
  AOI21X1 U31 ( .A0(n29), .A1(n101), .B0(sum[35]), .Y(n102) );
  INVX2 U32 ( .A(sum[1]), .Y(n2) );
  INVX2 U33 ( .A(sum[6]), .Y(n7) );
  INVX2 U34 ( .A(sum[3]), .Y(n4) );
  AOI21X1 U35 ( .A0(n127), .A1(n120), .B0(sum[39]), .Y(length[1]) );
  OAI211X1 U36 ( .A0(n119), .A1(n118), .B0(n30), .C0(n31), .Y(n120) );
  NAND2X1 U37 ( .A(n28), .B(n29), .Y(n118) );
  AOI31X1 U38 ( .A0(n6), .A1(n7), .A2(n105), .B0(n104), .Y(n107) );
  OR2X1 U39 ( .A(sum[7]), .B(sum[8]), .Y(n104) );
  OAI211X1 U40 ( .A0(sum[1]), .A1(sum[2]), .B0(n4), .C0(n5), .Y(n105) );
  AOI31X1 U41 ( .A0(n12), .A1(n13), .A2(n109), .B0(n108), .Y(n111) );
  OR2X1 U42 ( .A(sum[15]), .B(sum[16]), .Y(n108) );
  OAI211X1 U43 ( .A0(n107), .A1(n106), .B0(n10), .C0(n11), .Y(n109) );
  NAND2X1 U44 ( .A(n9), .B(n8), .Y(n106) );
  AOI31X1 U45 ( .A0(n18), .A1(n19), .A2(n113), .B0(n112), .Y(n115) );
  OR2X1 U46 ( .A(sum[23]), .B(sum[24]), .Y(n112) );
  OAI211X1 U47 ( .A0(n111), .A1(n110), .B0(n16), .C0(n17), .Y(n113) );
  INVX2 U48 ( .A(sum[20]), .Y(n17) );
  AOI31X1 U49 ( .A0(n26), .A1(n27), .A2(n117), .B0(n116), .Y(n119) );
  OR2X1 U50 ( .A(sum[31]), .B(sum[32]), .Y(n116) );
  OAI211X1 U51 ( .A0(n115), .A1(n114), .B0(n24), .C0(n25), .Y(n117) );
  NAND2X1 U52 ( .A(n22), .B(n23), .Y(n114) );
  INVX2 U53 ( .A(sum[5]), .Y(n6) );
  INVX2 U54 ( .A(sum[4]), .Y(n5) );
  INVX2 U55 ( .A(sum[10]), .Y(n9) );
  INVX2 U56 ( .A(sum[9]), .Y(n8) );
  INVX2 U57 ( .A(sum[11]), .Y(n10) );
  INVX2 U58 ( .A(sum[14]), .Y(n13) );
  INVX2 U59 ( .A(sum[12]), .Y(n11) );
  INVX2 U60 ( .A(sum[13]), .Y(n12) );
  INVX2 U61 ( .A(sum[18]), .Y(n15) );
  INVX2 U62 ( .A(sum[17]), .Y(n14) );
  INVX2 U63 ( .A(sum[19]), .Y(n16) );
  NOR3X1 U64 ( .A(sum[7]), .B(sum[9]), .C(sum[8]), .Y(n121) );
  AOI2BB1X1 U65 ( .A0N(n128), .A1N(n136), .B0(sum[39]), .Y(length[2]) );
  NOR2X1 U66 ( .A(n126), .B(n135), .Y(n128) );
  AOI31X1 U67 ( .A0(n125), .A1(n20), .A2(n124), .B0(n131), .Y(n126) );
  INVX2 U68 ( .A(sum[22]), .Y(n19) );
  INVX2 U69 ( .A(sum[21]), .Y(n18) );
  NAND4BBX1 U70 ( .AN(n130), .BN(sum[7]), .C(n9), .D(n129), .Y(n133) );
  NOR2X1 U71 ( .A(sum[9]), .B(sum[8]), .Y(n129) );
  OAI31X1 U72 ( .A0(n135), .A1(n134), .A2(n136), .B0(n1), .Y(length[3]) );
  INVX2 U73 ( .A(sum[39]), .Y(n1) );
  AOI31X1 U74 ( .A0(n138), .A1(n133), .A2(n137), .B0(n21), .Y(n134) );
  NOR4BX1 U75 ( .AN(n132), .B(n131), .C(sum[23]), .D(sum[24]), .Y(n139) );
  NOR2X1 U76 ( .A(sum[26]), .B(sum[25]), .Y(n132) );
  INVX2 U77 ( .A(sum[30]), .Y(n27) );
  INVX2 U78 ( .A(sum[26]), .Y(n23) );
  INVX2 U79 ( .A(sum[27]), .Y(n24) );
  INVX2 U80 ( .A(sum[25]), .Y(n22) );
  NOR4X1 U81 ( .A(sum[19]), .B(sum[20]), .C(sum[21]), .D(sum[22]), .Y(n138) );
  OR4X2 U82 ( .A(sum[31]), .B(sum[32]), .C(sum[33]), .D(sum[34]), .Y(n135) );
  OR3X2 U83 ( .A(n136), .B(sum[39]), .C(n135), .Y(length[5]) );
  NOR4X1 U84 ( .A(sum[15]), .B(sum[16]), .C(sum[17]), .D(sum[18]), .Y(n137) );
  INVX2 U85 ( .A(sum[28]), .Y(n25) );
  INVX2 U86 ( .A(sum[29]), .Y(n26) );
  NOR3X1 U87 ( .A(sum[24]), .B(sum[26]), .C(sum[25]), .Y(n124) );
  INVX2 U88 ( .A(sum[23]), .Y(n20) );
  NOR2X1 U89 ( .A(sum[38]), .B(sum[37]), .Y(n127) );
  INVX2 U90 ( .A(sum[35]), .Y(n30) );
  INVX2 U91 ( .A(sum[33]), .Y(n28) );
  INVX2 U92 ( .A(sum[34]), .Y(n29) );
  INVX2 U93 ( .A(sum[36]), .Y(n31) );
endmodule


module compare_8 ( clk, rst, sum, length );
  input [39:0] sum;
  output [5:0] length;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139;

  NAND2X1 U3 ( .A(n14), .B(n15), .Y(n110) );
  OAI2BB1X1 U4 ( .A0N(n3), .A1N(n137), .B0(n138), .Y(n125) );
  INVX2 U5 ( .A(n123), .Y(n3) );
  AOI31X1 U6 ( .A0(n122), .A1(n9), .A2(n121), .B0(n130), .Y(n123) );
  NAND4X1 U7 ( .A(n4), .B(n5), .C(n6), .D(n7), .Y(n122) );
  NAND4X1 U8 ( .A(n10), .B(n11), .C(n12), .D(n13), .Y(n130) );
  NAND4X1 U9 ( .A(n24), .B(n25), .C(n26), .D(n27), .Y(n131) );
  INVX2 U10 ( .A(n139), .Y(n21) );
  AOI31X1 U11 ( .A0(n139), .A1(n138), .A2(n137), .B0(length[5]), .Y(length[4])
         );
  NAND3X1 U12 ( .A(n30), .B(n31), .C(n127), .Y(n136) );
  OAI21X1 U13 ( .A0(n96), .A1(sum[24]), .B0(n22), .Y(n97) );
  AOI21X1 U14 ( .A0(n19), .A1(n95), .B0(sum[23]), .Y(n96) );
  OAI21X1 U15 ( .A0(n94), .A1(sum[20]), .B0(n18), .Y(n95) );
  AOI21X1 U16 ( .A0(n15), .A1(n93), .B0(sum[19]), .Y(n94) );
  OAI21X1 U17 ( .A0(n92), .A1(sum[16]), .B0(n14), .Y(n93) );
  AOI21X1 U18 ( .A0(n13), .A1(n91), .B0(sum[15]), .Y(n92) );
  OAI21X1 U19 ( .A0(n90), .A1(sum[12]), .B0(n12), .Y(n91) );
  AOI21X1 U20 ( .A0(n9), .A1(n89), .B0(sum[11]), .Y(n90) );
  OAI21X1 U21 ( .A0(n88), .A1(sum[8]), .B0(n8), .Y(n89) );
  AOI21X1 U22 ( .A0(n7), .A1(n87), .B0(sum[7]), .Y(n88) );
  OAI21X1 U23 ( .A0(n86), .A1(sum[4]), .B0(n6), .Y(n87) );
  AOI2BB1X1 U24 ( .A0N(n2), .A1N(sum[2]), .B0(sum[3]), .Y(n86) );
  OAI21X1 U25 ( .A0(n100), .A1(sum[32]), .B0(n28), .Y(n101) );
  AOI21X1 U26 ( .A0(n27), .A1(n99), .B0(sum[31]), .Y(n100) );
  OAI21X1 U27 ( .A0(n98), .A1(sum[28]), .B0(n26), .Y(n99) );
  AOI21X1 U28 ( .A0(n23), .A1(n97), .B0(sum[27]), .Y(n98) );
  AOI2BB1X1 U29 ( .A0N(sum[38]), .A1N(n103), .B0(sum[39]), .Y(length[0]) );
  AOI2BB1X1 U30 ( .A0N(n102), .A1N(sum[36]), .B0(sum[37]), .Y(n103) );
  AOI21X1 U31 ( .A0(n29), .A1(n101), .B0(sum[35]), .Y(n102) );
  INVX2 U32 ( .A(sum[1]), .Y(n2) );
  INVX2 U33 ( .A(sum[6]), .Y(n7) );
  INVX2 U34 ( .A(sum[3]), .Y(n4) );
  AOI21X1 U35 ( .A0(n127), .A1(n120), .B0(sum[39]), .Y(length[1]) );
  OAI211X1 U36 ( .A0(n119), .A1(n118), .B0(n30), .C0(n31), .Y(n120) );
  NAND2X1 U37 ( .A(n28), .B(n29), .Y(n118) );
  AOI31X1 U38 ( .A0(n6), .A1(n7), .A2(n105), .B0(n104), .Y(n107) );
  OR2X1 U39 ( .A(sum[7]), .B(sum[8]), .Y(n104) );
  OAI211X1 U40 ( .A0(sum[1]), .A1(sum[2]), .B0(n4), .C0(n5), .Y(n105) );
  AOI31X1 U41 ( .A0(n12), .A1(n13), .A2(n109), .B0(n108), .Y(n111) );
  OR2X1 U42 ( .A(sum[15]), .B(sum[16]), .Y(n108) );
  OAI211X1 U43 ( .A0(n107), .A1(n106), .B0(n10), .C0(n11), .Y(n109) );
  NAND2X1 U44 ( .A(n9), .B(n8), .Y(n106) );
  AOI31X1 U45 ( .A0(n18), .A1(n19), .A2(n113), .B0(n112), .Y(n115) );
  OR2X1 U46 ( .A(sum[23]), .B(sum[24]), .Y(n112) );
  OAI211X1 U47 ( .A0(n111), .A1(n110), .B0(n16), .C0(n17), .Y(n113) );
  INVX2 U48 ( .A(sum[20]), .Y(n17) );
  AOI31X1 U49 ( .A0(n26), .A1(n27), .A2(n117), .B0(n116), .Y(n119) );
  OR2X1 U50 ( .A(sum[31]), .B(sum[32]), .Y(n116) );
  OAI211X1 U51 ( .A0(n115), .A1(n114), .B0(n24), .C0(n25), .Y(n117) );
  NAND2X1 U52 ( .A(n22), .B(n23), .Y(n114) );
  INVX2 U53 ( .A(sum[5]), .Y(n6) );
  INVX2 U54 ( .A(sum[4]), .Y(n5) );
  INVX2 U55 ( .A(sum[10]), .Y(n9) );
  INVX2 U56 ( .A(sum[9]), .Y(n8) );
  INVX2 U57 ( .A(sum[11]), .Y(n10) );
  INVX2 U58 ( .A(sum[14]), .Y(n13) );
  INVX2 U59 ( .A(sum[13]), .Y(n12) );
  INVX2 U60 ( .A(sum[12]), .Y(n11) );
  INVX2 U61 ( .A(sum[18]), .Y(n15) );
  INVX2 U62 ( .A(sum[17]), .Y(n14) );
  INVX2 U63 ( .A(sum[19]), .Y(n16) );
  NOR3X1 U64 ( .A(sum[7]), .B(sum[9]), .C(sum[8]), .Y(n121) );
  AOI2BB1X1 U65 ( .A0N(n128), .A1N(n136), .B0(sum[39]), .Y(length[2]) );
  NOR2X1 U66 ( .A(n126), .B(n135), .Y(n128) );
  AOI31X1 U67 ( .A0(n125), .A1(n20), .A2(n124), .B0(n131), .Y(n126) );
  INVX2 U68 ( .A(sum[22]), .Y(n19) );
  INVX2 U69 ( .A(sum[21]), .Y(n18) );
  NAND4BBX1 U70 ( .AN(n130), .BN(sum[7]), .C(n9), .D(n129), .Y(n133) );
  NOR2X1 U71 ( .A(sum[9]), .B(sum[8]), .Y(n129) );
  OAI31X1 U72 ( .A0(n135), .A1(n134), .A2(n136), .B0(n1), .Y(length[3]) );
  INVX2 U73 ( .A(sum[39]), .Y(n1) );
  AOI31X1 U74 ( .A0(n138), .A1(n133), .A2(n137), .B0(n21), .Y(n134) );
  INVX2 U75 ( .A(sum[26]), .Y(n23) );
  INVX2 U76 ( .A(sum[25]), .Y(n22) );
  NOR4BX1 U77 ( .AN(n132), .B(n131), .C(sum[23]), .D(sum[24]), .Y(n139) );
  NOR2X1 U78 ( .A(sum[26]), .B(sum[25]), .Y(n132) );
  INVX2 U79 ( .A(sum[30]), .Y(n27) );
  INVX2 U80 ( .A(sum[27]), .Y(n24) );
  OR4X2 U81 ( .A(sum[31]), .B(sum[32]), .C(sum[33]), .D(sum[34]), .Y(n135) );
  OR3X2 U82 ( .A(n136), .B(sum[39]), .C(n135), .Y(length[5]) );
  NOR4X1 U83 ( .A(sum[19]), .B(sum[20]), .C(sum[21]), .D(sum[22]), .Y(n138) );
  NOR4X1 U84 ( .A(sum[15]), .B(sum[16]), .C(sum[17]), .D(sum[18]), .Y(n137) );
  INVX2 U85 ( .A(sum[29]), .Y(n26) );
  INVX2 U86 ( .A(sum[28]), .Y(n25) );
  NOR3X1 U87 ( .A(sum[24]), .B(sum[26]), .C(sum[25]), .Y(n124) );
  INVX2 U88 ( .A(sum[23]), .Y(n20) );
  NOR2X1 U89 ( .A(sum[38]), .B(sum[37]), .Y(n127) );
  INVX2 U90 ( .A(sum[35]), .Y(n30) );
  INVX2 U91 ( .A(sum[33]), .Y(n28) );
  INVX2 U92 ( .A(sum[34]), .Y(n29) );
  INVX2 U93 ( .A(sum[36]), .Y(n31) );
endmodule


module compare_9 ( clk, rst, sum, length );
  input [39:0] sum;
  output [5:0] length;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139;

  NAND2X1 U3 ( .A(n14), .B(n15), .Y(n110) );
  OAI2BB1X1 U4 ( .A0N(n3), .A1N(n137), .B0(n138), .Y(n125) );
  INVX2 U5 ( .A(n123), .Y(n3) );
  AOI31X1 U6 ( .A0(n122), .A1(n9), .A2(n121), .B0(n130), .Y(n123) );
  NAND4X1 U7 ( .A(n4), .B(n5), .C(n6), .D(n7), .Y(n122) );
  NAND4X1 U8 ( .A(n10), .B(n11), .C(n12), .D(n13), .Y(n130) );
  NAND4X1 U9 ( .A(n24), .B(n25), .C(n26), .D(n27), .Y(n131) );
  INVX2 U10 ( .A(n139), .Y(n21) );
  AOI31X1 U11 ( .A0(n139), .A1(n138), .A2(n137), .B0(length[5]), .Y(length[4])
         );
  NAND3X1 U12 ( .A(n30), .B(n31), .C(n127), .Y(n136) );
  OAI21X1 U13 ( .A0(n88), .A1(sum[8]), .B0(n8), .Y(n89) );
  AOI21X1 U14 ( .A0(n7), .A1(n87), .B0(sum[7]), .Y(n88) );
  OAI21X1 U15 ( .A0(n86), .A1(sum[4]), .B0(n6), .Y(n87) );
  AOI2BB1X1 U16 ( .A0N(n2), .A1N(sum[2]), .B0(sum[3]), .Y(n86) );
  OAI21X1 U17 ( .A0(n96), .A1(sum[24]), .B0(n22), .Y(n97) );
  AOI21X1 U18 ( .A0(n19), .A1(n95), .B0(sum[23]), .Y(n96) );
  OAI21X1 U19 ( .A0(n94), .A1(sum[20]), .B0(n18), .Y(n95) );
  AOI21X1 U20 ( .A0(n15), .A1(n93), .B0(sum[19]), .Y(n94) );
  OAI21X1 U21 ( .A0(n92), .A1(sum[16]), .B0(n14), .Y(n93) );
  AOI21X1 U22 ( .A0(n13), .A1(n91), .B0(sum[15]), .Y(n92) );
  OAI21X1 U23 ( .A0(n90), .A1(sum[12]), .B0(n12), .Y(n91) );
  AOI21X1 U24 ( .A0(n9), .A1(n89), .B0(sum[11]), .Y(n90) );
  OAI21X1 U25 ( .A0(n100), .A1(sum[32]), .B0(n28), .Y(n101) );
  AOI21X1 U26 ( .A0(n27), .A1(n99), .B0(sum[31]), .Y(n100) );
  OAI21X1 U27 ( .A0(n98), .A1(sum[28]), .B0(n26), .Y(n99) );
  AOI21X1 U28 ( .A0(n23), .A1(n97), .B0(sum[27]), .Y(n98) );
  INVX2 U29 ( .A(sum[1]), .Y(n2) );
  AOI2BB1X1 U30 ( .A0N(sum[38]), .A1N(n103), .B0(sum[39]), .Y(length[0]) );
  AOI2BB1X1 U31 ( .A0N(n102), .A1N(sum[36]), .B0(sum[37]), .Y(n103) );
  AOI21X1 U32 ( .A0(n29), .A1(n101), .B0(sum[35]), .Y(n102) );
  INVX2 U33 ( .A(sum[5]), .Y(n6) );
  INVX2 U34 ( .A(sum[6]), .Y(n7) );
  INVX2 U35 ( .A(sum[3]), .Y(n4) );
  AOI21X1 U36 ( .A0(n127), .A1(n120), .B0(sum[39]), .Y(length[1]) );
  OAI211X1 U37 ( .A0(n119), .A1(n118), .B0(n30), .C0(n31), .Y(n120) );
  NAND2X1 U38 ( .A(n28), .B(n29), .Y(n118) );
  AOI31X1 U39 ( .A0(n6), .A1(n7), .A2(n105), .B0(n104), .Y(n107) );
  OR2X1 U40 ( .A(sum[7]), .B(sum[8]), .Y(n104) );
  OAI211X1 U41 ( .A0(sum[1]), .A1(sum[2]), .B0(n4), .C0(n5), .Y(n105) );
  AOI31X1 U42 ( .A0(n12), .A1(n13), .A2(n109), .B0(n108), .Y(n111) );
  OR2X1 U43 ( .A(sum[15]), .B(sum[16]), .Y(n108) );
  OAI211X1 U44 ( .A0(n107), .A1(n106), .B0(n10), .C0(n11), .Y(n109) );
  NAND2X1 U45 ( .A(n9), .B(n8), .Y(n106) );
  AOI31X1 U46 ( .A0(n18), .A1(n19), .A2(n113), .B0(n112), .Y(n115) );
  OR2X1 U47 ( .A(sum[23]), .B(sum[24]), .Y(n112) );
  OAI211X1 U48 ( .A0(n111), .A1(n110), .B0(n16), .C0(n17), .Y(n113) );
  INVX2 U49 ( .A(sum[19]), .Y(n16) );
  AOI31X1 U50 ( .A0(n26), .A1(n27), .A2(n117), .B0(n116), .Y(n119) );
  OR2X1 U51 ( .A(sum[31]), .B(sum[32]), .Y(n116) );
  OAI211X1 U52 ( .A0(n115), .A1(n114), .B0(n24), .C0(n25), .Y(n117) );
  NAND2X1 U53 ( .A(n22), .B(n23), .Y(n114) );
  INVX2 U54 ( .A(sum[4]), .Y(n5) );
  INVX2 U55 ( .A(sum[9]), .Y(n8) );
  INVX2 U56 ( .A(sum[10]), .Y(n9) );
  INVX2 U57 ( .A(sum[13]), .Y(n12) );
  INVX2 U58 ( .A(sum[14]), .Y(n13) );
  INVX2 U59 ( .A(sum[12]), .Y(n11) );
  INVX2 U60 ( .A(sum[11]), .Y(n10) );
  INVX2 U61 ( .A(sum[17]), .Y(n14) );
  INVX2 U62 ( .A(sum[18]), .Y(n15) );
  INVX2 U63 ( .A(sum[21]), .Y(n18) );
  INVX2 U64 ( .A(sum[20]), .Y(n17) );
  NOR3X1 U65 ( .A(sum[7]), .B(sum[9]), .C(sum[8]), .Y(n121) );
  AOI2BB1X1 U66 ( .A0N(n128), .A1N(n136), .B0(sum[39]), .Y(length[2]) );
  NOR2X1 U67 ( .A(n126), .B(n135), .Y(n128) );
  AOI31X1 U68 ( .A0(n125), .A1(n20), .A2(n124), .B0(n131), .Y(n126) );
  INVX2 U69 ( .A(sum[22]), .Y(n19) );
  INVX2 U70 ( .A(sum[25]), .Y(n22) );
  INVX2 U71 ( .A(sum[26]), .Y(n23) );
  NAND4BBX1 U72 ( .AN(n130), .BN(sum[7]), .C(n9), .D(n129), .Y(n133) );
  NOR2X1 U73 ( .A(sum[9]), .B(sum[8]), .Y(n129) );
  OAI31X1 U74 ( .A0(n135), .A1(n134), .A2(n136), .B0(n1), .Y(length[3]) );
  INVX2 U75 ( .A(sum[39]), .Y(n1) );
  AOI31X1 U76 ( .A0(n138), .A1(n133), .A2(n137), .B0(n21), .Y(n134) );
  NOR4BX1 U77 ( .AN(n132), .B(n131), .C(sum[23]), .D(sum[24]), .Y(n139) );
  NOR2X1 U78 ( .A(sum[26]), .B(sum[25]), .Y(n132) );
  INVX2 U79 ( .A(sum[28]), .Y(n25) );
  INVX2 U80 ( .A(sum[27]), .Y(n24) );
  INVX2 U81 ( .A(sum[30]), .Y(n27) );
  INVX2 U82 ( .A(sum[29]), .Y(n26) );
  OR4X2 U83 ( .A(sum[31]), .B(sum[32]), .C(sum[33]), .D(sum[34]), .Y(n135) );
  OR3X2 U84 ( .A(n136), .B(sum[39]), .C(n135), .Y(length[5]) );
  NOR4X1 U85 ( .A(sum[19]), .B(sum[20]), .C(sum[21]), .D(sum[22]), .Y(n138) );
  NOR4X1 U86 ( .A(sum[15]), .B(sum[16]), .C(sum[17]), .D(sum[18]), .Y(n137) );
  NOR3X1 U87 ( .A(sum[24]), .B(sum[26]), .C(sum[25]), .Y(n124) );
  INVX2 U88 ( .A(sum[23]), .Y(n20) );
  INVX2 U89 ( .A(sum[33]), .Y(n28) );
  NOR2X1 U90 ( .A(sum[38]), .B(sum[37]), .Y(n127) );
  INVX2 U91 ( .A(sum[36]), .Y(n31) );
  INVX2 U92 ( .A(sum[35]), .Y(n30) );
  INVX2 U93 ( .A(sum[34]), .Y(n29) );
endmodule


module compare_10 ( clk, rst, sum, length );
  input [39:0] sum;
  output [5:0] length;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139;

  NAND2X1 U3 ( .A(n14), .B(n15), .Y(n110) );
  OAI2BB1X1 U4 ( .A0N(n3), .A1N(n137), .B0(n138), .Y(n125) );
  INVX2 U5 ( .A(n123), .Y(n3) );
  AOI31X1 U6 ( .A0(n122), .A1(n9), .A2(n121), .B0(n130), .Y(n123) );
  NAND4X1 U7 ( .A(n4), .B(n5), .C(n6), .D(n7), .Y(n122) );
  NAND4X1 U8 ( .A(n10), .B(n11), .C(n12), .D(n13), .Y(n130) );
  INVX2 U9 ( .A(n139), .Y(n21) );
  NAND4X1 U10 ( .A(n24), .B(n25), .C(n26), .D(n27), .Y(n131) );
  AOI31X1 U11 ( .A0(n139), .A1(n138), .A2(n137), .B0(length[5]), .Y(length[4])
         );
  NAND3X1 U12 ( .A(n30), .B(n31), .C(n127), .Y(n136) );
  OAI21X1 U13 ( .A0(n96), .A1(sum[24]), .B0(n22), .Y(n97) );
  AOI21X1 U14 ( .A0(n19), .A1(n95), .B0(sum[23]), .Y(n96) );
  OAI21X1 U15 ( .A0(n94), .A1(sum[20]), .B0(n18), .Y(n95) );
  AOI21X1 U16 ( .A0(n15), .A1(n93), .B0(sum[19]), .Y(n94) );
  OAI21X1 U17 ( .A0(n88), .A1(sum[8]), .B0(n8), .Y(n89) );
  AOI21X1 U18 ( .A0(n7), .A1(n87), .B0(sum[7]), .Y(n88) );
  OAI21X1 U19 ( .A0(n86), .A1(sum[4]), .B0(n6), .Y(n87) );
  AOI2BB1X1 U20 ( .A0N(n2), .A1N(sum[2]), .B0(sum[3]), .Y(n86) );
  OAI21X1 U21 ( .A0(n100), .A1(sum[32]), .B0(n28), .Y(n101) );
  AOI21X1 U22 ( .A0(n27), .A1(n99), .B0(sum[31]), .Y(n100) );
  OAI21X1 U23 ( .A0(n98), .A1(sum[28]), .B0(n26), .Y(n99) );
  AOI21X1 U24 ( .A0(n23), .A1(n97), .B0(sum[27]), .Y(n98) );
  OAI21X1 U25 ( .A0(n92), .A1(sum[16]), .B0(n14), .Y(n93) );
  AOI21X1 U26 ( .A0(n13), .A1(n91), .B0(sum[15]), .Y(n92) );
  OAI21X1 U27 ( .A0(n90), .A1(sum[12]), .B0(n12), .Y(n91) );
  AOI21X1 U28 ( .A0(n9), .A1(n89), .B0(sum[11]), .Y(n90) );
  INVX2 U29 ( .A(sum[1]), .Y(n2) );
  AOI2BB1X1 U30 ( .A0N(sum[38]), .A1N(n103), .B0(sum[39]), .Y(length[0]) );
  AOI2BB1X1 U31 ( .A0N(n102), .A1N(sum[36]), .B0(sum[37]), .Y(n103) );
  AOI21X1 U32 ( .A0(n29), .A1(n101), .B0(sum[35]), .Y(n102) );
  INVX2 U33 ( .A(sum[5]), .Y(n6) );
  INVX2 U34 ( .A(sum[4]), .Y(n5) );
  AOI21X1 U35 ( .A0(n127), .A1(n120), .B0(sum[39]), .Y(length[1]) );
  OAI211X1 U36 ( .A0(n119), .A1(n118), .B0(n30), .C0(n31), .Y(n120) );
  NAND2X1 U37 ( .A(n28), .B(n29), .Y(n118) );
  AOI31X1 U38 ( .A0(n6), .A1(n7), .A2(n105), .B0(n104), .Y(n107) );
  OR2X1 U39 ( .A(sum[7]), .B(sum[8]), .Y(n104) );
  OAI211X1 U40 ( .A0(sum[1]), .A1(sum[2]), .B0(n4), .C0(n5), .Y(n105) );
  AOI31X1 U41 ( .A0(n12), .A1(n13), .A2(n109), .B0(n108), .Y(n111) );
  OR2X1 U42 ( .A(sum[15]), .B(sum[16]), .Y(n108) );
  OAI211X1 U43 ( .A0(n107), .A1(n106), .B0(n10), .C0(n11), .Y(n109) );
  NAND2X1 U44 ( .A(n9), .B(n8), .Y(n106) );
  AOI31X1 U45 ( .A0(n18), .A1(n19), .A2(n113), .B0(n112), .Y(n115) );
  OR2X1 U46 ( .A(sum[23]), .B(sum[24]), .Y(n112) );
  OAI211X1 U47 ( .A0(n111), .A1(n110), .B0(n16), .C0(n17), .Y(n113) );
  INVX2 U48 ( .A(sum[19]), .Y(n16) );
  AOI31X1 U49 ( .A0(n26), .A1(n27), .A2(n117), .B0(n116), .Y(n119) );
  OR2X1 U50 ( .A(sum[31]), .B(sum[32]), .Y(n116) );
  OAI211X1 U51 ( .A0(n115), .A1(n114), .B0(n24), .C0(n25), .Y(n117) );
  NAND2X1 U52 ( .A(n22), .B(n23), .Y(n114) );
  INVX2 U53 ( .A(sum[3]), .Y(n4) );
  INVX2 U54 ( .A(sum[6]), .Y(n7) );
  INVX2 U55 ( .A(sum[9]), .Y(n8) );
  INVX2 U56 ( .A(sum[10]), .Y(n9) );
  INVX2 U57 ( .A(sum[13]), .Y(n12) );
  INVX2 U58 ( .A(sum[12]), .Y(n11) );
  INVX2 U59 ( .A(sum[11]), .Y(n10) );
  INVX2 U60 ( .A(sum[14]), .Y(n13) );
  INVX2 U61 ( .A(sum[17]), .Y(n14) );
  INVX2 U62 ( .A(sum[18]), .Y(n15) );
  INVX2 U63 ( .A(sum[21]), .Y(n18) );
  INVX2 U64 ( .A(sum[20]), .Y(n17) );
  NOR3X1 U65 ( .A(sum[7]), .B(sum[9]), .C(sum[8]), .Y(n121) );
  AOI2BB1X1 U66 ( .A0N(n128), .A1N(n136), .B0(sum[39]), .Y(length[2]) );
  NOR2X1 U67 ( .A(n126), .B(n135), .Y(n128) );
  AOI31X1 U68 ( .A0(n125), .A1(n20), .A2(n124), .B0(n131), .Y(n126) );
  INVX2 U69 ( .A(sum[22]), .Y(n19) );
  INVX2 U70 ( .A(sum[25]), .Y(n22) );
  NAND4BBX1 U71 ( .AN(n130), .BN(sum[7]), .C(n9), .D(n129), .Y(n133) );
  NOR2X1 U72 ( .A(sum[9]), .B(sum[8]), .Y(n129) );
  OAI31X1 U73 ( .A0(n135), .A1(n134), .A2(n136), .B0(n1), .Y(length[3]) );
  INVX2 U74 ( .A(sum[39]), .Y(n1) );
  AOI31X1 U75 ( .A0(n138), .A1(n133), .A2(n137), .B0(n21), .Y(n134) );
  NOR4BX1 U76 ( .AN(n132), .B(n131), .C(sum[23]), .D(sum[24]), .Y(n139) );
  NOR2X1 U77 ( .A(sum[26]), .B(sum[25]), .Y(n132) );
  INVX2 U78 ( .A(sum[28]), .Y(n25) );
  INVX2 U79 ( .A(sum[26]), .Y(n23) );
  INVX2 U80 ( .A(sum[30]), .Y(n27) );
  INVX2 U81 ( .A(sum[27]), .Y(n24) );
  INVX2 U82 ( .A(sum[29]), .Y(n26) );
  OR4X2 U83 ( .A(sum[31]), .B(sum[32]), .C(sum[33]), .D(sum[34]), .Y(n135) );
  OR3X2 U84 ( .A(n136), .B(sum[39]), .C(n135), .Y(length[5]) );
  NOR4X1 U85 ( .A(sum[15]), .B(sum[16]), .C(sum[17]), .D(sum[18]), .Y(n137) );
  NOR4X1 U86 ( .A(sum[19]), .B(sum[20]), .C(sum[21]), .D(sum[22]), .Y(n138) );
  NOR3X1 U87 ( .A(sum[24]), .B(sum[26]), .C(sum[25]), .Y(n124) );
  INVX2 U88 ( .A(sum[23]), .Y(n20) );
  NOR2X1 U89 ( .A(sum[38]), .B(sum[37]), .Y(n127) );
  INVX2 U90 ( .A(sum[33]), .Y(n28) );
  INVX2 U91 ( .A(sum[36]), .Y(n31) );
  INVX2 U92 ( .A(sum[35]), .Y(n30) );
  INVX2 U93 ( .A(sum[34]), .Y(n29) );
endmodule


module compare_11 ( clk, rst, sum, length );
  input [39:0] sum;
  output [5:0] length;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139;

  NAND2X1 U3 ( .A(n14), .B(n15), .Y(n110) );
  OAI2BB1X1 U4 ( .A0N(n3), .A1N(n137), .B0(n138), .Y(n125) );
  INVX2 U5 ( .A(n123), .Y(n3) );
  AOI31X1 U6 ( .A0(n122), .A1(n9), .A2(n121), .B0(n130), .Y(n123) );
  NAND4X1 U7 ( .A(n4), .B(n5), .C(n6), .D(n7), .Y(n122) );
  NAND4X1 U8 ( .A(n10), .B(n11), .C(n12), .D(n13), .Y(n130) );
  NAND4X1 U9 ( .A(n24), .B(n25), .C(n26), .D(n27), .Y(n131) );
  INVX2 U10 ( .A(n139), .Y(n21) );
  AOI31X1 U11 ( .A0(n139), .A1(n138), .A2(n137), .B0(length[5]), .Y(length[4])
         );
  NAND3X1 U12 ( .A(n30), .B(n31), .C(n127), .Y(n136) );
  OAI21X1 U13 ( .A0(n96), .A1(sum[24]), .B0(n22), .Y(n97) );
  AOI21X1 U14 ( .A0(n19), .A1(n95), .B0(sum[23]), .Y(n96) );
  OAI21X1 U15 ( .A0(n94), .A1(sum[20]), .B0(n18), .Y(n95) );
  AOI21X1 U16 ( .A0(n15), .A1(n93), .B0(sum[19]), .Y(n94) );
  OAI21X1 U17 ( .A0(n92), .A1(sum[16]), .B0(n14), .Y(n93) );
  AOI21X1 U18 ( .A0(n13), .A1(n91), .B0(sum[15]), .Y(n92) );
  OAI21X1 U19 ( .A0(n90), .A1(sum[12]), .B0(n12), .Y(n91) );
  AOI21X1 U20 ( .A0(n9), .A1(n89), .B0(sum[11]), .Y(n90) );
  OAI21X1 U21 ( .A0(n100), .A1(sum[32]), .B0(n28), .Y(n101) );
  AOI21X1 U22 ( .A0(n27), .A1(n99), .B0(sum[31]), .Y(n100) );
  OAI21X1 U23 ( .A0(n98), .A1(sum[28]), .B0(n26), .Y(n99) );
  AOI21X1 U24 ( .A0(n23), .A1(n97), .B0(sum[27]), .Y(n98) );
  OAI21X1 U25 ( .A0(n88), .A1(sum[8]), .B0(n8), .Y(n89) );
  AOI21X1 U26 ( .A0(n7), .A1(n87), .B0(sum[7]), .Y(n88) );
  OAI21X1 U27 ( .A0(n86), .A1(sum[4]), .B0(n6), .Y(n87) );
  AOI2BB1X1 U28 ( .A0N(n2), .A1N(sum[2]), .B0(sum[3]), .Y(n86) );
  INVX2 U29 ( .A(sum[1]), .Y(n2) );
  AOI2BB1X1 U30 ( .A0N(sum[38]), .A1N(n103), .B0(sum[39]), .Y(length[0]) );
  AOI2BB1X1 U31 ( .A0N(n102), .A1N(sum[36]), .B0(sum[37]), .Y(n103) );
  AOI21X1 U32 ( .A0(n29), .A1(n101), .B0(sum[35]), .Y(n102) );
  INVX2 U33 ( .A(sum[5]), .Y(n6) );
  INVX2 U34 ( .A(sum[6]), .Y(n7) );
  INVX2 U35 ( .A(sum[3]), .Y(n4) );
  AOI21X1 U36 ( .A0(n127), .A1(n120), .B0(sum[39]), .Y(length[1]) );
  OAI211X1 U37 ( .A0(n119), .A1(n118), .B0(n30), .C0(n31), .Y(n120) );
  NAND2X1 U38 ( .A(n28), .B(n29), .Y(n118) );
  AOI31X1 U39 ( .A0(n6), .A1(n7), .A2(n105), .B0(n104), .Y(n107) );
  OR2X1 U40 ( .A(sum[7]), .B(sum[8]), .Y(n104) );
  OAI211X1 U41 ( .A0(sum[1]), .A1(sum[2]), .B0(n4), .C0(n5), .Y(n105) );
  AOI31X1 U42 ( .A0(n12), .A1(n13), .A2(n109), .B0(n108), .Y(n111) );
  OR2X1 U43 ( .A(sum[15]), .B(sum[16]), .Y(n108) );
  OAI211X1 U44 ( .A0(n107), .A1(n106), .B0(n10), .C0(n11), .Y(n109) );
  NAND2X1 U45 ( .A(n9), .B(n8), .Y(n106) );
  AOI31X1 U46 ( .A0(n18), .A1(n19), .A2(n113), .B0(n112), .Y(n115) );
  OR2X1 U47 ( .A(sum[23]), .B(sum[24]), .Y(n112) );
  OAI211X1 U48 ( .A0(n111), .A1(n110), .B0(n16), .C0(n17), .Y(n113) );
  INVX2 U49 ( .A(sum[19]), .Y(n16) );
  AOI31X1 U50 ( .A0(n26), .A1(n27), .A2(n117), .B0(n116), .Y(n119) );
  OR2X1 U51 ( .A(sum[31]), .B(sum[32]), .Y(n116) );
  OAI211X1 U52 ( .A0(n115), .A1(n114), .B0(n24), .C0(n25), .Y(n117) );
  NAND2X1 U53 ( .A(n22), .B(n23), .Y(n114) );
  INVX2 U54 ( .A(sum[9]), .Y(n8) );
  INVX2 U55 ( .A(sum[4]), .Y(n5) );
  INVX2 U56 ( .A(sum[10]), .Y(n9) );
  INVX2 U57 ( .A(sum[13]), .Y(n12) );
  INVX2 U58 ( .A(sum[14]), .Y(n13) );
  INVX2 U59 ( .A(sum[12]), .Y(n11) );
  INVX2 U60 ( .A(sum[11]), .Y(n10) );
  INVX2 U61 ( .A(sum[17]), .Y(n14) );
  INVX2 U62 ( .A(sum[18]), .Y(n15) );
  INVX2 U63 ( .A(sum[21]), .Y(n18) );
  INVX2 U64 ( .A(sum[20]), .Y(n17) );
  NOR3X1 U65 ( .A(sum[7]), .B(sum[9]), .C(sum[8]), .Y(n121) );
  AOI2BB1X1 U66 ( .A0N(n128), .A1N(n136), .B0(sum[39]), .Y(length[2]) );
  NOR2X1 U67 ( .A(n126), .B(n135), .Y(n128) );
  AOI31X1 U68 ( .A0(n125), .A1(n20), .A2(n124), .B0(n131), .Y(n126) );
  INVX2 U69 ( .A(sum[22]), .Y(n19) );
  INVX2 U70 ( .A(sum[25]), .Y(n22) );
  INVX2 U71 ( .A(sum[26]), .Y(n23) );
  NAND4BBX1 U72 ( .AN(n130), .BN(sum[7]), .C(n9), .D(n129), .Y(n133) );
  NOR2X1 U73 ( .A(sum[9]), .B(sum[8]), .Y(n129) );
  OAI31X1 U74 ( .A0(n135), .A1(n134), .A2(n136), .B0(n1), .Y(length[3]) );
  INVX2 U75 ( .A(sum[39]), .Y(n1) );
  AOI31X1 U76 ( .A0(n138), .A1(n133), .A2(n137), .B0(n21), .Y(n134) );
  NOR4BX1 U77 ( .AN(n132), .B(n131), .C(sum[23]), .D(sum[24]), .Y(n139) );
  NOR2X1 U78 ( .A(sum[26]), .B(sum[25]), .Y(n132) );
  INVX2 U79 ( .A(sum[28]), .Y(n25) );
  INVX2 U80 ( .A(sum[30]), .Y(n27) );
  INVX2 U81 ( .A(sum[27]), .Y(n24) );
  INVX2 U82 ( .A(sum[29]), .Y(n26) );
  OR4X2 U83 ( .A(sum[31]), .B(sum[32]), .C(sum[33]), .D(sum[34]), .Y(n135) );
  OR3X2 U84 ( .A(n136), .B(sum[39]), .C(n135), .Y(length[5]) );
  NOR4X1 U85 ( .A(sum[19]), .B(sum[20]), .C(sum[21]), .D(sum[22]), .Y(n138) );
  NOR4X1 U86 ( .A(sum[15]), .B(sum[16]), .C(sum[17]), .D(sum[18]), .Y(n137) );
  NOR3X1 U87 ( .A(sum[24]), .B(sum[26]), .C(sum[25]), .Y(n124) );
  INVX2 U88 ( .A(sum[23]), .Y(n20) );
  NOR2X1 U89 ( .A(sum[38]), .B(sum[37]), .Y(n127) );
  INVX2 U90 ( .A(sum[33]), .Y(n28) );
  INVX2 U91 ( .A(sum[36]), .Y(n31) );
  INVX2 U92 ( .A(sum[35]), .Y(n30) );
  INVX2 U93 ( .A(sum[34]), .Y(n29) );
endmodule


module compare_12 ( clk, rst, sum, length );
  input [39:0] sum;
  output [5:0] length;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139;

  NAND2X1 U3 ( .A(n14), .B(n15), .Y(n110) );
  OAI2BB1X1 U4 ( .A0N(n3), .A1N(n137), .B0(n138), .Y(n125) );
  INVX2 U5 ( .A(n123), .Y(n3) );
  AOI31X1 U6 ( .A0(n122), .A1(n9), .A2(n121), .B0(n130), .Y(n123) );
  NAND4X1 U7 ( .A(n4), .B(n5), .C(n6), .D(n7), .Y(n122) );
  NAND4X1 U8 ( .A(n10), .B(n11), .C(n12), .D(n13), .Y(n130) );
  NAND4X1 U9 ( .A(n24), .B(n25), .C(n26), .D(n27), .Y(n131) );
  INVX2 U10 ( .A(n139), .Y(n21) );
  AOI31X1 U11 ( .A0(n139), .A1(n138), .A2(n137), .B0(length[5]), .Y(length[4])
         );
  NAND3X1 U12 ( .A(n30), .B(n31), .C(n127), .Y(n136) );
  OAI21X1 U13 ( .A0(n88), .A1(sum[8]), .B0(n8), .Y(n89) );
  AOI21X1 U14 ( .A0(n7), .A1(n87), .B0(sum[7]), .Y(n88) );
  OAI21X1 U15 ( .A0(n86), .A1(sum[4]), .B0(n6), .Y(n87) );
  AOI2BB1X1 U16 ( .A0N(n2), .A1N(sum[2]), .B0(sum[3]), .Y(n86) );
  OAI21X1 U17 ( .A0(n96), .A1(sum[24]), .B0(n22), .Y(n97) );
  AOI21X1 U18 ( .A0(n19), .A1(n95), .B0(sum[23]), .Y(n96) );
  OAI21X1 U19 ( .A0(n94), .A1(sum[20]), .B0(n18), .Y(n95) );
  AOI21X1 U20 ( .A0(n15), .A1(n93), .B0(sum[19]), .Y(n94) );
  OAI21X1 U21 ( .A0(n92), .A1(sum[16]), .B0(n14), .Y(n93) );
  AOI21X1 U22 ( .A0(n13), .A1(n91), .B0(sum[15]), .Y(n92) );
  OAI21X1 U23 ( .A0(n90), .A1(sum[12]), .B0(n12), .Y(n91) );
  AOI21X1 U24 ( .A0(n9), .A1(n89), .B0(sum[11]), .Y(n90) );
  OAI21X1 U25 ( .A0(n100), .A1(sum[32]), .B0(n28), .Y(n101) );
  AOI21X1 U26 ( .A0(n27), .A1(n99), .B0(sum[31]), .Y(n100) );
  OAI21X1 U27 ( .A0(n98), .A1(sum[28]), .B0(n26), .Y(n99) );
  AOI21X1 U28 ( .A0(n23), .A1(n97), .B0(sum[27]), .Y(n98) );
  INVX2 U29 ( .A(sum[1]), .Y(n2) );
  AOI2BB1X1 U30 ( .A0N(sum[38]), .A1N(n103), .B0(sum[39]), .Y(length[0]) );
  AOI2BB1X1 U31 ( .A0N(n102), .A1N(sum[36]), .B0(sum[37]), .Y(n103) );
  AOI21X1 U32 ( .A0(n29), .A1(n101), .B0(sum[35]), .Y(n102) );
  INVX2 U33 ( .A(sum[5]), .Y(n6) );
  INVX2 U34 ( .A(sum[6]), .Y(n7) );
  INVX2 U35 ( .A(sum[4]), .Y(n5) );
  AOI21X1 U36 ( .A0(n127), .A1(n120), .B0(sum[39]), .Y(length[1]) );
  OAI211X1 U37 ( .A0(n119), .A1(n118), .B0(n30), .C0(n31), .Y(n120) );
  NAND2X1 U38 ( .A(n28), .B(n29), .Y(n118) );
  AOI31X1 U39 ( .A0(n6), .A1(n7), .A2(n105), .B0(n104), .Y(n107) );
  OR2X1 U40 ( .A(sum[7]), .B(sum[8]), .Y(n104) );
  OAI211X1 U41 ( .A0(sum[1]), .A1(sum[2]), .B0(n4), .C0(n5), .Y(n105) );
  AOI31X1 U42 ( .A0(n12), .A1(n13), .A2(n109), .B0(n108), .Y(n111) );
  OR2X1 U43 ( .A(sum[15]), .B(sum[16]), .Y(n108) );
  OAI211X1 U44 ( .A0(n107), .A1(n106), .B0(n10), .C0(n11), .Y(n109) );
  NAND2X1 U45 ( .A(n9), .B(n8), .Y(n106) );
  AOI31X1 U46 ( .A0(n18), .A1(n19), .A2(n113), .B0(n112), .Y(n115) );
  OR2X1 U47 ( .A(sum[23]), .B(sum[24]), .Y(n112) );
  OAI211X1 U48 ( .A0(n111), .A1(n110), .B0(n16), .C0(n17), .Y(n113) );
  INVX2 U49 ( .A(sum[19]), .Y(n16) );
  AOI31X1 U50 ( .A0(n26), .A1(n27), .A2(n117), .B0(n116), .Y(n119) );
  OR2X1 U51 ( .A(sum[31]), .B(sum[32]), .Y(n116) );
  OAI211X1 U52 ( .A0(n115), .A1(n114), .B0(n24), .C0(n25), .Y(n117) );
  NAND2X1 U53 ( .A(n22), .B(n23), .Y(n114) );
  INVX2 U54 ( .A(sum[3]), .Y(n4) );
  INVX2 U55 ( .A(sum[9]), .Y(n8) );
  INVX2 U56 ( .A(sum[10]), .Y(n9) );
  INVX2 U57 ( .A(sum[13]), .Y(n12) );
  INVX2 U58 ( .A(sum[14]), .Y(n13) );
  INVX2 U59 ( .A(sum[12]), .Y(n11) );
  INVX2 U60 ( .A(sum[11]), .Y(n10) );
  INVX2 U61 ( .A(sum[17]), .Y(n14) );
  INVX2 U62 ( .A(sum[18]), .Y(n15) );
  INVX2 U63 ( .A(sum[21]), .Y(n18) );
  INVX2 U64 ( .A(sum[20]), .Y(n17) );
  NOR3X1 U65 ( .A(sum[7]), .B(sum[9]), .C(sum[8]), .Y(n121) );
  AOI2BB1X1 U66 ( .A0N(n128), .A1N(n136), .B0(sum[39]), .Y(length[2]) );
  NOR2X1 U67 ( .A(n126), .B(n135), .Y(n128) );
  AOI31X1 U68 ( .A0(n125), .A1(n20), .A2(n124), .B0(n131), .Y(n126) );
  INVX2 U69 ( .A(sum[22]), .Y(n19) );
  INVX2 U70 ( .A(sum[25]), .Y(n22) );
  INVX2 U71 ( .A(sum[26]), .Y(n23) );
  NAND4BBX1 U72 ( .AN(n130), .BN(sum[7]), .C(n9), .D(n129), .Y(n133) );
  NOR2X1 U73 ( .A(sum[9]), .B(sum[8]), .Y(n129) );
  OAI31X1 U74 ( .A0(n135), .A1(n134), .A2(n136), .B0(n1), .Y(length[3]) );
  INVX2 U75 ( .A(sum[39]), .Y(n1) );
  AOI31X1 U76 ( .A0(n138), .A1(n133), .A2(n137), .B0(n21), .Y(n134) );
  NOR4BX1 U77 ( .AN(n132), .B(n131), .C(sum[23]), .D(sum[24]), .Y(n139) );
  NOR2X1 U78 ( .A(sum[26]), .B(sum[25]), .Y(n132) );
  INVX2 U79 ( .A(sum[28]), .Y(n25) );
  INVX2 U80 ( .A(sum[29]), .Y(n26) );
  INVX2 U81 ( .A(sum[30]), .Y(n27) );
  INVX2 U82 ( .A(sum[27]), .Y(n24) );
  OR4X2 U83 ( .A(sum[31]), .B(sum[32]), .C(sum[33]), .D(sum[34]), .Y(n135) );
  OR3X2 U84 ( .A(n136), .B(sum[39]), .C(n135), .Y(length[5]) );
  NOR4X1 U85 ( .A(sum[19]), .B(sum[20]), .C(sum[21]), .D(sum[22]), .Y(n138) );
  NOR4X1 U86 ( .A(sum[15]), .B(sum[16]), .C(sum[17]), .D(sum[18]), .Y(n137) );
  NOR3X1 U87 ( .A(sum[24]), .B(sum[26]), .C(sum[25]), .Y(n124) );
  INVX2 U88 ( .A(sum[23]), .Y(n20) );
  NOR2X1 U89 ( .A(sum[38]), .B(sum[37]), .Y(n127) );
  INVX2 U90 ( .A(sum[33]), .Y(n28) );
  INVX2 U91 ( .A(sum[36]), .Y(n31) );
  INVX2 U92 ( .A(sum[35]), .Y(n30) );
  INVX2 U93 ( .A(sum[34]), .Y(n29) );
endmodule


module compare_13 ( clk, rst, sum, length );
  input [39:0] sum;
  output [5:0] length;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139;

  NAND2X1 U3 ( .A(n14), .B(n15), .Y(n110) );
  OAI2BB1X1 U4 ( .A0N(n3), .A1N(n137), .B0(n138), .Y(n125) );
  INVX2 U5 ( .A(n123), .Y(n3) );
  AOI31X1 U6 ( .A0(n122), .A1(n9), .A2(n121), .B0(n130), .Y(n123) );
  NAND4X1 U7 ( .A(n4), .B(n5), .C(n6), .D(n7), .Y(n122) );
  NAND4X1 U8 ( .A(n10), .B(n11), .C(n12), .D(n13), .Y(n130) );
  INVX2 U9 ( .A(n139), .Y(n21) );
  NAND4X1 U10 ( .A(n24), .B(n25), .C(n26), .D(n27), .Y(n131) );
  AOI31X1 U11 ( .A0(n139), .A1(n138), .A2(n137), .B0(length[5]), .Y(length[4])
         );
  NAND3X1 U12 ( .A(n30), .B(n31), .C(n127), .Y(n136) );
  OAI21X1 U13 ( .A0(n96), .A1(sum[24]), .B0(n22), .Y(n97) );
  AOI21X1 U14 ( .A0(n19), .A1(n95), .B0(sum[23]), .Y(n96) );
  OAI21X1 U15 ( .A0(n94), .A1(sum[20]), .B0(n18), .Y(n95) );
  AOI21X1 U16 ( .A0(n15), .A1(n93), .B0(sum[19]), .Y(n94) );
  OAI21X1 U17 ( .A0(n88), .A1(sum[8]), .B0(n8), .Y(n89) );
  AOI21X1 U18 ( .A0(n7), .A1(n87), .B0(sum[7]), .Y(n88) );
  OAI21X1 U19 ( .A0(n86), .A1(sum[4]), .B0(n6), .Y(n87) );
  AOI2BB1X1 U20 ( .A0N(n2), .A1N(sum[2]), .B0(sum[3]), .Y(n86) );
  OAI21X1 U21 ( .A0(n92), .A1(sum[16]), .B0(n14), .Y(n93) );
  AOI21X1 U22 ( .A0(n13), .A1(n91), .B0(sum[15]), .Y(n92) );
  OAI21X1 U23 ( .A0(n90), .A1(sum[12]), .B0(n12), .Y(n91) );
  AOI21X1 U24 ( .A0(n9), .A1(n89), .B0(sum[11]), .Y(n90) );
  OAI21X1 U25 ( .A0(n100), .A1(sum[32]), .B0(n28), .Y(n101) );
  AOI21X1 U26 ( .A0(n27), .A1(n99), .B0(sum[31]), .Y(n100) );
  OAI21X1 U27 ( .A0(n98), .A1(sum[28]), .B0(n26), .Y(n99) );
  AOI21X1 U28 ( .A0(n23), .A1(n97), .B0(sum[27]), .Y(n98) );
  INVX2 U29 ( .A(sum[1]), .Y(n2) );
  AOI2BB1X1 U30 ( .A0N(sum[38]), .A1N(n103), .B0(sum[39]), .Y(length[0]) );
  AOI2BB1X1 U31 ( .A0N(n102), .A1N(sum[36]), .B0(sum[37]), .Y(n103) );
  AOI21X1 U32 ( .A0(n29), .A1(n101), .B0(sum[35]), .Y(n102) );
  INVX2 U33 ( .A(sum[5]), .Y(n6) );
  INVX2 U34 ( .A(sum[6]), .Y(n7) );
  AOI31X1 U35 ( .A0(n12), .A1(n13), .A2(n109), .B0(n108), .Y(n111) );
  OR2X1 U36 ( .A(sum[15]), .B(sum[16]), .Y(n108) );
  OAI211X1 U37 ( .A0(n107), .A1(n106), .B0(n10), .C0(n11), .Y(n109) );
  NAND2X1 U38 ( .A(n9), .B(n8), .Y(n106) );
  INVX2 U39 ( .A(sum[4]), .Y(n5) );
  AOI21X1 U40 ( .A0(n127), .A1(n120), .B0(sum[39]), .Y(length[1]) );
  OAI211X1 U41 ( .A0(n119), .A1(n118), .B0(n30), .C0(n31), .Y(n120) );
  NAND2X1 U42 ( .A(n28), .B(n29), .Y(n118) );
  AOI31X1 U43 ( .A0(n6), .A1(n7), .A2(n105), .B0(n104), .Y(n107) );
  OR2X1 U44 ( .A(sum[7]), .B(sum[8]), .Y(n104) );
  OAI211X1 U45 ( .A0(sum[1]), .A1(sum[2]), .B0(n4), .C0(n5), .Y(n105) );
  AOI31X1 U46 ( .A0(n18), .A1(n19), .A2(n113), .B0(n112), .Y(n115) );
  OR2X1 U47 ( .A(sum[23]), .B(sum[24]), .Y(n112) );
  OAI211X1 U48 ( .A0(n111), .A1(n110), .B0(n16), .C0(n17), .Y(n113) );
  INVX2 U49 ( .A(sum[19]), .Y(n16) );
  AOI31X1 U50 ( .A0(n26), .A1(n27), .A2(n117), .B0(n116), .Y(n119) );
  OR2X1 U51 ( .A(sum[31]), .B(sum[32]), .Y(n116) );
  OAI211X1 U52 ( .A0(n115), .A1(n114), .B0(n24), .C0(n25), .Y(n117) );
  NAND2X1 U53 ( .A(n22), .B(n23), .Y(n114) );
  INVX2 U54 ( .A(sum[3]), .Y(n4) );
  INVX2 U55 ( .A(sum[9]), .Y(n8) );
  INVX2 U56 ( .A(sum[10]), .Y(n9) );
  INVX2 U57 ( .A(sum[13]), .Y(n12) );
  INVX2 U58 ( .A(sum[14]), .Y(n13) );
  INVX2 U59 ( .A(sum[12]), .Y(n11) );
  INVX2 U60 ( .A(sum[11]), .Y(n10) );
  INVX2 U61 ( .A(sum[17]), .Y(n14) );
  INVX2 U62 ( .A(sum[18]), .Y(n15) );
  INVX2 U63 ( .A(sum[21]), .Y(n18) );
  INVX2 U64 ( .A(sum[20]), .Y(n17) );
  NOR3X1 U65 ( .A(sum[7]), .B(sum[9]), .C(sum[8]), .Y(n121) );
  AOI2BB1X1 U66 ( .A0N(n128), .A1N(n136), .B0(sum[39]), .Y(length[2]) );
  NOR2X1 U67 ( .A(n126), .B(n135), .Y(n128) );
  AOI31X1 U68 ( .A0(n125), .A1(n20), .A2(n124), .B0(n131), .Y(n126) );
  INVX2 U69 ( .A(sum[22]), .Y(n19) );
  INVX2 U70 ( .A(sum[25]), .Y(n22) );
  INVX2 U71 ( .A(sum[26]), .Y(n23) );
  NAND4BBX1 U72 ( .AN(n130), .BN(sum[7]), .C(n9), .D(n129), .Y(n133) );
  NOR2X1 U73 ( .A(sum[9]), .B(sum[8]), .Y(n129) );
  OAI31X1 U74 ( .A0(n135), .A1(n134), .A2(n136), .B0(n1), .Y(length[3]) );
  INVX2 U75 ( .A(sum[39]), .Y(n1) );
  AOI31X1 U76 ( .A0(n138), .A1(n133), .A2(n137), .B0(n21), .Y(n134) );
  NOR4BX1 U77 ( .AN(n132), .B(n131), .C(sum[23]), .D(sum[24]), .Y(n139) );
  NOR2X1 U78 ( .A(sum[26]), .B(sum[25]), .Y(n132) );
  INVX2 U79 ( .A(sum[28]), .Y(n25) );
  INVX2 U80 ( .A(sum[30]), .Y(n27) );
  INVX2 U81 ( .A(sum[27]), .Y(n24) );
  INVX2 U82 ( .A(sum[29]), .Y(n26) );
  OR4X2 U83 ( .A(sum[31]), .B(sum[32]), .C(sum[33]), .D(sum[34]), .Y(n135) );
  OR3X2 U84 ( .A(n136), .B(sum[39]), .C(n135), .Y(length[5]) );
  NOR4X1 U85 ( .A(sum[19]), .B(sum[20]), .C(sum[21]), .D(sum[22]), .Y(n138) );
  NOR4X1 U86 ( .A(sum[15]), .B(sum[16]), .C(sum[17]), .D(sum[18]), .Y(n137) );
  NOR3X1 U87 ( .A(sum[24]), .B(sum[26]), .C(sum[25]), .Y(n124) );
  INVX2 U88 ( .A(sum[23]), .Y(n20) );
  NOR2X1 U89 ( .A(sum[38]), .B(sum[37]), .Y(n127) );
  INVX2 U90 ( .A(sum[33]), .Y(n28) );
  INVX2 U91 ( .A(sum[36]), .Y(n31) );
  INVX2 U92 ( .A(sum[35]), .Y(n30) );
  INVX2 U93 ( .A(sum[34]), .Y(n29) );
endmodule


module compare_0 ( clk, rst, sum, length );
  input [39:0] sum;
  output [5:0] length;
  input clk, rst;
  wire   n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31;

  NAND2X1 U3 ( .A(n14), .B(n15), .Y(n61) );
  OAI2BB1X1 U4 ( .A0N(n3), .A1N(n34), .B0(n33), .Y(n46) );
  INVX2 U5 ( .A(n48), .Y(n3) );
  AOI31X1 U6 ( .A0(n49), .A1(n9), .A2(n50), .B0(n41), .Y(n48) );
  NAND4X1 U7 ( .A(n4), .B(n5), .C(n6), .D(n7), .Y(n49) );
  NAND4X1 U8 ( .A(n10), .B(n11), .C(n12), .D(n13), .Y(n41) );
  NAND4X1 U9 ( .A(n24), .B(n25), .C(n26), .D(n27), .Y(n40) );
  INVX2 U10 ( .A(n32), .Y(n21) );
  AOI31X1 U11 ( .A0(n32), .A1(n33), .A2(n34), .B0(length[5]), .Y(length[4]) );
  NAND3X1 U12 ( .A(n30), .B(n31), .C(n44), .Y(n35) );
  OAI21X1 U13 ( .A0(n75), .A1(sum[24]), .B0(n22), .Y(n74) );
  AOI21X1 U14 ( .A0(n19), .A1(n76), .B0(sum[23]), .Y(n75) );
  OAI21X1 U15 ( .A0(n77), .A1(sum[20]), .B0(n18), .Y(n76) );
  AOI21X1 U16 ( .A0(n15), .A1(n78), .B0(sum[19]), .Y(n77) );
  OAI21X1 U17 ( .A0(n83), .A1(sum[8]), .B0(n8), .Y(n82) );
  AOI21X1 U18 ( .A0(n7), .A1(n84), .B0(sum[7]), .Y(n83) );
  OAI21X1 U19 ( .A0(n85), .A1(sum[4]), .B0(n6), .Y(n84) );
  AOI2BB1X1 U20 ( .A0N(n2), .A1N(sum[2]), .B0(sum[3]), .Y(n85) );
  OAI21X1 U21 ( .A0(n71), .A1(sum[32]), .B0(n28), .Y(n70) );
  AOI21X1 U22 ( .A0(n27), .A1(n72), .B0(sum[31]), .Y(n71) );
  OAI21X1 U23 ( .A0(n73), .A1(sum[28]), .B0(n26), .Y(n72) );
  AOI21X1 U24 ( .A0(n23), .A1(n74), .B0(sum[27]), .Y(n73) );
  OAI21X1 U25 ( .A0(n79), .A1(sum[16]), .B0(n14), .Y(n78) );
  AOI21X1 U26 ( .A0(n13), .A1(n80), .B0(sum[15]), .Y(n79) );
  OAI21X1 U27 ( .A0(n81), .A1(sum[12]), .B0(n12), .Y(n80) );
  AOI21X1 U28 ( .A0(n9), .A1(n82), .B0(sum[11]), .Y(n81) );
  INVX2 U29 ( .A(sum[1]), .Y(n2) );
  AOI2BB1X1 U30 ( .A0N(sum[38]), .A1N(n68), .B0(sum[39]), .Y(length[0]) );
  AOI2BB1X1 U31 ( .A0N(n69), .A1N(sum[36]), .B0(sum[37]), .Y(n68) );
  AOI21X1 U32 ( .A0(n29), .A1(n70), .B0(sum[35]), .Y(n69) );
  INVX2 U33 ( .A(sum[5]), .Y(n6) );
  INVX2 U34 ( .A(sum[6]), .Y(n7) );
  AOI31X1 U35 ( .A0(n18), .A1(n19), .A2(n58), .B0(n59), .Y(n56) );
  OR2X1 U36 ( .A(sum[23]), .B(sum[24]), .Y(n59) );
  OAI211X1 U37 ( .A0(n60), .A1(n61), .B0(n16), .C0(n17), .Y(n58) );
  INVX2 U38 ( .A(sum[19]), .Y(n16) );
  INVX2 U39 ( .A(sum[4]), .Y(n5) );
  AOI21X1 U40 ( .A0(n44), .A1(n51), .B0(sum[39]), .Y(length[1]) );
  OAI211X1 U41 ( .A0(n52), .A1(n53), .B0(n30), .C0(n31), .Y(n51) );
  NAND2X1 U42 ( .A(n28), .B(n29), .Y(n53) );
  AOI31X1 U43 ( .A0(n6), .A1(n7), .A2(n66), .B0(n67), .Y(n64) );
  OR2X1 U44 ( .A(sum[7]), .B(sum[8]), .Y(n67) );
  OAI211X1 U45 ( .A0(sum[1]), .A1(sum[2]), .B0(n4), .C0(n5), .Y(n66) );
  AOI31X1 U46 ( .A0(n12), .A1(n13), .A2(n62), .B0(n63), .Y(n60) );
  OR2X1 U47 ( .A(sum[15]), .B(sum[16]), .Y(n63) );
  OAI211X1 U48 ( .A0(n64), .A1(n65), .B0(n10), .C0(n11), .Y(n62) );
  NAND2X1 U49 ( .A(n9), .B(n8), .Y(n65) );
  AOI31X1 U50 ( .A0(n26), .A1(n27), .A2(n54), .B0(n55), .Y(n52) );
  OR2X1 U51 ( .A(sum[31]), .B(sum[32]), .Y(n55) );
  OAI211X1 U52 ( .A0(n56), .A1(n57), .B0(n24), .C0(n25), .Y(n54) );
  NAND2X1 U53 ( .A(n22), .B(n23), .Y(n57) );
  INVX2 U54 ( .A(sum[3]), .Y(n4) );
  INVX2 U55 ( .A(sum[9]), .Y(n8) );
  INVX2 U56 ( .A(sum[10]), .Y(n9) );
  INVX2 U57 ( .A(sum[13]), .Y(n12) );
  INVX2 U58 ( .A(sum[14]), .Y(n13) );
  INVX2 U59 ( .A(sum[12]), .Y(n11) );
  INVX2 U60 ( .A(sum[11]), .Y(n10) );
  INVX2 U61 ( .A(sum[17]), .Y(n14) );
  INVX2 U62 ( .A(sum[18]), .Y(n15) );
  INVX2 U63 ( .A(sum[21]), .Y(n18) );
  INVX2 U64 ( .A(sum[20]), .Y(n17) );
  NOR3X1 U65 ( .A(sum[7]), .B(sum[9]), .C(sum[8]), .Y(n50) );
  AOI2BB1X1 U66 ( .A0N(n43), .A1N(n35), .B0(sum[39]), .Y(length[2]) );
  NOR2X1 U67 ( .A(n45), .B(n36), .Y(n43) );
  AOI31X1 U68 ( .A0(n46), .A1(n20), .A2(n47), .B0(n40), .Y(n45) );
  INVX2 U69 ( .A(sum[22]), .Y(n19) );
  INVX2 U70 ( .A(sum[25]), .Y(n22) );
  INVX2 U71 ( .A(sum[26]), .Y(n23) );
  NAND4BBX1 U72 ( .AN(n41), .BN(sum[7]), .C(n9), .D(n42), .Y(n38) );
  NOR2X1 U73 ( .A(sum[9]), .B(sum[8]), .Y(n42) );
  OAI31X1 U74 ( .A0(n36), .A1(n37), .A2(n35), .B0(n1), .Y(length[3]) );
  INVX2 U75 ( .A(sum[39]), .Y(n1) );
  AOI31X1 U76 ( .A0(n33), .A1(n38), .A2(n34), .B0(n21), .Y(n37) );
  NOR4BX1 U77 ( .AN(n39), .B(n40), .C(sum[23]), .D(sum[24]), .Y(n32) );
  NOR2X1 U78 ( .A(sum[26]), .B(sum[25]), .Y(n39) );
  INVX2 U79 ( .A(sum[28]), .Y(n25) );
  INVX2 U80 ( .A(sum[29]), .Y(n26) );
  INVX2 U81 ( .A(sum[27]), .Y(n24) );
  INVX2 U82 ( .A(sum[30]), .Y(n27) );
  OR4X2 U83 ( .A(sum[31]), .B(sum[32]), .C(sum[33]), .D(sum[34]), .Y(n36) );
  OR3X2 U84 ( .A(n35), .B(sum[39]), .C(n36), .Y(length[5]) );
  NOR4X1 U85 ( .A(sum[19]), .B(sum[20]), .C(sum[21]), .D(sum[22]), .Y(n33) );
  NOR4X1 U86 ( .A(sum[15]), .B(sum[16]), .C(sum[17]), .D(sum[18]), .Y(n34) );
  NOR3X1 U87 ( .A(sum[24]), .B(sum[26]), .C(sum[25]), .Y(n47) );
  INVX2 U88 ( .A(sum[23]), .Y(n20) );
  NOR2X1 U89 ( .A(sum[38]), .B(sum[37]), .Y(n44) );
  INVX2 U90 ( .A(sum[33]), .Y(n28) );
  INVX2 U91 ( .A(sum[36]), .Y(n31) );
  INVX2 U92 ( .A(sum[35]), .Y(n30) );
  INVX2 U93 ( .A(sum[34]), .Y(n29) );
endmodule

